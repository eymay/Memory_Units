module Regfile (clk,
    rst,
    we0,
    rd_addr0,
    rd_addr1,
    rd_dout0,
    rd_dout1,
    wr_addr0,
    wr_din0);
 input clk;
 input rst;
 input we0;
 input [4:0] rd_addr0;
 input [4:0] rd_addr1;
 output [31:0] rd_dout0;
 output [31:0] rd_dout1;
 input [4:0] wr_addr0;
 input [31:0] wr_din0;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[16][0] ;
 wire \mem[16][10] ;
 wire \mem[16][11] ;
 wire \mem[16][12] ;
 wire \mem[16][13] ;
 wire \mem[16][14] ;
 wire \mem[16][15] ;
 wire \mem[16][16] ;
 wire \mem[16][17] ;
 wire \mem[16][18] ;
 wire \mem[16][19] ;
 wire \mem[16][1] ;
 wire \mem[16][20] ;
 wire \mem[16][21] ;
 wire \mem[16][22] ;
 wire \mem[16][23] ;
 wire \mem[16][24] ;
 wire \mem[16][25] ;
 wire \mem[16][26] ;
 wire \mem[16][27] ;
 wire \mem[16][28] ;
 wire \mem[16][29] ;
 wire \mem[16][2] ;
 wire \mem[16][30] ;
 wire \mem[16][31] ;
 wire \mem[16][3] ;
 wire \mem[16][4] ;
 wire \mem[16][5] ;
 wire \mem[16][6] ;
 wire \mem[16][7] ;
 wire \mem[16][8] ;
 wire \mem[16][9] ;
 wire \mem[17][0] ;
 wire \mem[17][10] ;
 wire \mem[17][11] ;
 wire \mem[17][12] ;
 wire \mem[17][13] ;
 wire \mem[17][14] ;
 wire \mem[17][15] ;
 wire \mem[17][16] ;
 wire \mem[17][17] ;
 wire \mem[17][18] ;
 wire \mem[17][19] ;
 wire \mem[17][1] ;
 wire \mem[17][20] ;
 wire \mem[17][21] ;
 wire \mem[17][22] ;
 wire \mem[17][23] ;
 wire \mem[17][24] ;
 wire \mem[17][25] ;
 wire \mem[17][26] ;
 wire \mem[17][27] ;
 wire \mem[17][28] ;
 wire \mem[17][29] ;
 wire \mem[17][2] ;
 wire \mem[17][30] ;
 wire \mem[17][31] ;
 wire \mem[17][3] ;
 wire \mem[17][4] ;
 wire \mem[17][5] ;
 wire \mem[17][6] ;
 wire \mem[17][7] ;
 wire \mem[17][8] ;
 wire \mem[17][9] ;
 wire \mem[18][0] ;
 wire \mem[18][10] ;
 wire \mem[18][11] ;
 wire \mem[18][12] ;
 wire \mem[18][13] ;
 wire \mem[18][14] ;
 wire \mem[18][15] ;
 wire \mem[18][16] ;
 wire \mem[18][17] ;
 wire \mem[18][18] ;
 wire \mem[18][19] ;
 wire \mem[18][1] ;
 wire \mem[18][20] ;
 wire \mem[18][21] ;
 wire \mem[18][22] ;
 wire \mem[18][23] ;
 wire \mem[18][24] ;
 wire \mem[18][25] ;
 wire \mem[18][26] ;
 wire \mem[18][27] ;
 wire \mem[18][28] ;
 wire \mem[18][29] ;
 wire \mem[18][2] ;
 wire \mem[18][30] ;
 wire \mem[18][31] ;
 wire \mem[18][3] ;
 wire \mem[18][4] ;
 wire \mem[18][5] ;
 wire \mem[18][6] ;
 wire \mem[18][7] ;
 wire \mem[18][8] ;
 wire \mem[18][9] ;
 wire \mem[19][0] ;
 wire \mem[19][10] ;
 wire \mem[19][11] ;
 wire \mem[19][12] ;
 wire \mem[19][13] ;
 wire \mem[19][14] ;
 wire \mem[19][15] ;
 wire \mem[19][16] ;
 wire \mem[19][17] ;
 wire \mem[19][18] ;
 wire \mem[19][19] ;
 wire \mem[19][1] ;
 wire \mem[19][20] ;
 wire \mem[19][21] ;
 wire \mem[19][22] ;
 wire \mem[19][23] ;
 wire \mem[19][24] ;
 wire \mem[19][25] ;
 wire \mem[19][26] ;
 wire \mem[19][27] ;
 wire \mem[19][28] ;
 wire \mem[19][29] ;
 wire \mem[19][2] ;
 wire \mem[19][30] ;
 wire \mem[19][31] ;
 wire \mem[19][3] ;
 wire \mem[19][4] ;
 wire \mem[19][5] ;
 wire \mem[19][6] ;
 wire \mem[19][7] ;
 wire \mem[19][8] ;
 wire \mem[19][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[20][0] ;
 wire \mem[20][10] ;
 wire \mem[20][11] ;
 wire \mem[20][12] ;
 wire \mem[20][13] ;
 wire \mem[20][14] ;
 wire \mem[20][15] ;
 wire \mem[20][16] ;
 wire \mem[20][17] ;
 wire \mem[20][18] ;
 wire \mem[20][19] ;
 wire \mem[20][1] ;
 wire \mem[20][20] ;
 wire \mem[20][21] ;
 wire \mem[20][22] ;
 wire \mem[20][23] ;
 wire \mem[20][24] ;
 wire \mem[20][25] ;
 wire \mem[20][26] ;
 wire \mem[20][27] ;
 wire \mem[20][28] ;
 wire \mem[20][29] ;
 wire \mem[20][2] ;
 wire \mem[20][30] ;
 wire \mem[20][31] ;
 wire \mem[20][3] ;
 wire \mem[20][4] ;
 wire \mem[20][5] ;
 wire \mem[20][6] ;
 wire \mem[20][7] ;
 wire \mem[20][8] ;
 wire \mem[20][9] ;
 wire \mem[21][0] ;
 wire \mem[21][10] ;
 wire \mem[21][11] ;
 wire \mem[21][12] ;
 wire \mem[21][13] ;
 wire \mem[21][14] ;
 wire \mem[21][15] ;
 wire \mem[21][16] ;
 wire \mem[21][17] ;
 wire \mem[21][18] ;
 wire \mem[21][19] ;
 wire \mem[21][1] ;
 wire \mem[21][20] ;
 wire \mem[21][21] ;
 wire \mem[21][22] ;
 wire \mem[21][23] ;
 wire \mem[21][24] ;
 wire \mem[21][25] ;
 wire \mem[21][26] ;
 wire \mem[21][27] ;
 wire \mem[21][28] ;
 wire \mem[21][29] ;
 wire \mem[21][2] ;
 wire \mem[21][30] ;
 wire \mem[21][31] ;
 wire \mem[21][3] ;
 wire \mem[21][4] ;
 wire \mem[21][5] ;
 wire \mem[21][6] ;
 wire \mem[21][7] ;
 wire \mem[21][8] ;
 wire \mem[21][9] ;
 wire \mem[22][0] ;
 wire \mem[22][10] ;
 wire \mem[22][11] ;
 wire \mem[22][12] ;
 wire \mem[22][13] ;
 wire \mem[22][14] ;
 wire \mem[22][15] ;
 wire \mem[22][16] ;
 wire \mem[22][17] ;
 wire \mem[22][18] ;
 wire \mem[22][19] ;
 wire \mem[22][1] ;
 wire \mem[22][20] ;
 wire \mem[22][21] ;
 wire \mem[22][22] ;
 wire \mem[22][23] ;
 wire \mem[22][24] ;
 wire \mem[22][25] ;
 wire \mem[22][26] ;
 wire \mem[22][27] ;
 wire \mem[22][28] ;
 wire \mem[22][29] ;
 wire \mem[22][2] ;
 wire \mem[22][30] ;
 wire \mem[22][31] ;
 wire \mem[22][3] ;
 wire \mem[22][4] ;
 wire \mem[22][5] ;
 wire \mem[22][6] ;
 wire \mem[22][7] ;
 wire \mem[22][8] ;
 wire \mem[22][9] ;
 wire \mem[23][0] ;
 wire \mem[23][10] ;
 wire \mem[23][11] ;
 wire \mem[23][12] ;
 wire \mem[23][13] ;
 wire \mem[23][14] ;
 wire \mem[23][15] ;
 wire \mem[23][16] ;
 wire \mem[23][17] ;
 wire \mem[23][18] ;
 wire \mem[23][19] ;
 wire \mem[23][1] ;
 wire \mem[23][20] ;
 wire \mem[23][21] ;
 wire \mem[23][22] ;
 wire \mem[23][23] ;
 wire \mem[23][24] ;
 wire \mem[23][25] ;
 wire \mem[23][26] ;
 wire \mem[23][27] ;
 wire \mem[23][28] ;
 wire \mem[23][29] ;
 wire \mem[23][2] ;
 wire \mem[23][30] ;
 wire \mem[23][31] ;
 wire \mem[23][3] ;
 wire \mem[23][4] ;
 wire \mem[23][5] ;
 wire \mem[23][6] ;
 wire \mem[23][7] ;
 wire \mem[23][8] ;
 wire \mem[23][9] ;
 wire \mem[24][0] ;
 wire \mem[24][10] ;
 wire \mem[24][11] ;
 wire \mem[24][12] ;
 wire \mem[24][13] ;
 wire \mem[24][14] ;
 wire \mem[24][15] ;
 wire \mem[24][16] ;
 wire \mem[24][17] ;
 wire \mem[24][18] ;
 wire \mem[24][19] ;
 wire \mem[24][1] ;
 wire \mem[24][20] ;
 wire \mem[24][21] ;
 wire \mem[24][22] ;
 wire \mem[24][23] ;
 wire \mem[24][24] ;
 wire \mem[24][25] ;
 wire \mem[24][26] ;
 wire \mem[24][27] ;
 wire \mem[24][28] ;
 wire \mem[24][29] ;
 wire \mem[24][2] ;
 wire \mem[24][30] ;
 wire \mem[24][31] ;
 wire \mem[24][3] ;
 wire \mem[24][4] ;
 wire \mem[24][5] ;
 wire \mem[24][6] ;
 wire \mem[24][7] ;
 wire \mem[24][8] ;
 wire \mem[24][9] ;
 wire \mem[25][0] ;
 wire \mem[25][10] ;
 wire \mem[25][11] ;
 wire \mem[25][12] ;
 wire \mem[25][13] ;
 wire \mem[25][14] ;
 wire \mem[25][15] ;
 wire \mem[25][16] ;
 wire \mem[25][17] ;
 wire \mem[25][18] ;
 wire \mem[25][19] ;
 wire \mem[25][1] ;
 wire \mem[25][20] ;
 wire \mem[25][21] ;
 wire \mem[25][22] ;
 wire \mem[25][23] ;
 wire \mem[25][24] ;
 wire \mem[25][25] ;
 wire \mem[25][26] ;
 wire \mem[25][27] ;
 wire \mem[25][28] ;
 wire \mem[25][29] ;
 wire \mem[25][2] ;
 wire \mem[25][30] ;
 wire \mem[25][31] ;
 wire \mem[25][3] ;
 wire \mem[25][4] ;
 wire \mem[25][5] ;
 wire \mem[25][6] ;
 wire \mem[25][7] ;
 wire \mem[25][8] ;
 wire \mem[25][9] ;
 wire \mem[26][0] ;
 wire \mem[26][10] ;
 wire \mem[26][11] ;
 wire \mem[26][12] ;
 wire \mem[26][13] ;
 wire \mem[26][14] ;
 wire \mem[26][15] ;
 wire \mem[26][16] ;
 wire \mem[26][17] ;
 wire \mem[26][18] ;
 wire \mem[26][19] ;
 wire \mem[26][1] ;
 wire \mem[26][20] ;
 wire \mem[26][21] ;
 wire \mem[26][22] ;
 wire \mem[26][23] ;
 wire \mem[26][24] ;
 wire \mem[26][25] ;
 wire \mem[26][26] ;
 wire \mem[26][27] ;
 wire \mem[26][28] ;
 wire \mem[26][29] ;
 wire \mem[26][2] ;
 wire \mem[26][30] ;
 wire \mem[26][31] ;
 wire \mem[26][3] ;
 wire \mem[26][4] ;
 wire \mem[26][5] ;
 wire \mem[26][6] ;
 wire \mem[26][7] ;
 wire \mem[26][8] ;
 wire \mem[26][9] ;
 wire \mem[27][0] ;
 wire \mem[27][10] ;
 wire \mem[27][11] ;
 wire \mem[27][12] ;
 wire \mem[27][13] ;
 wire \mem[27][14] ;
 wire \mem[27][15] ;
 wire \mem[27][16] ;
 wire \mem[27][17] ;
 wire \mem[27][18] ;
 wire \mem[27][19] ;
 wire \mem[27][1] ;
 wire \mem[27][20] ;
 wire \mem[27][21] ;
 wire \mem[27][22] ;
 wire \mem[27][23] ;
 wire \mem[27][24] ;
 wire \mem[27][25] ;
 wire \mem[27][26] ;
 wire \mem[27][27] ;
 wire \mem[27][28] ;
 wire \mem[27][29] ;
 wire \mem[27][2] ;
 wire \mem[27][30] ;
 wire \mem[27][31] ;
 wire \mem[27][3] ;
 wire \mem[27][4] ;
 wire \mem[27][5] ;
 wire \mem[27][6] ;
 wire \mem[27][7] ;
 wire \mem[27][8] ;
 wire \mem[27][9] ;
 wire \mem[28][0] ;
 wire \mem[28][10] ;
 wire \mem[28][11] ;
 wire \mem[28][12] ;
 wire \mem[28][13] ;
 wire \mem[28][14] ;
 wire \mem[28][15] ;
 wire \mem[28][16] ;
 wire \mem[28][17] ;
 wire \mem[28][18] ;
 wire \mem[28][19] ;
 wire \mem[28][1] ;
 wire \mem[28][20] ;
 wire \mem[28][21] ;
 wire \mem[28][22] ;
 wire \mem[28][23] ;
 wire \mem[28][24] ;
 wire \mem[28][25] ;
 wire \mem[28][26] ;
 wire \mem[28][27] ;
 wire \mem[28][28] ;
 wire \mem[28][29] ;
 wire \mem[28][2] ;
 wire \mem[28][30] ;
 wire \mem[28][31] ;
 wire \mem[28][3] ;
 wire \mem[28][4] ;
 wire \mem[28][5] ;
 wire \mem[28][6] ;
 wire \mem[28][7] ;
 wire \mem[28][8] ;
 wire \mem[28][9] ;
 wire \mem[29][0] ;
 wire \mem[29][10] ;
 wire \mem[29][11] ;
 wire \mem[29][12] ;
 wire \mem[29][13] ;
 wire \mem[29][14] ;
 wire \mem[29][15] ;
 wire \mem[29][16] ;
 wire \mem[29][17] ;
 wire \mem[29][18] ;
 wire \mem[29][19] ;
 wire \mem[29][1] ;
 wire \mem[29][20] ;
 wire \mem[29][21] ;
 wire \mem[29][22] ;
 wire \mem[29][23] ;
 wire \mem[29][24] ;
 wire \mem[29][25] ;
 wire \mem[29][26] ;
 wire \mem[29][27] ;
 wire \mem[29][28] ;
 wire \mem[29][29] ;
 wire \mem[29][2] ;
 wire \mem[29][30] ;
 wire \mem[29][31] ;
 wire \mem[29][3] ;
 wire \mem[29][4] ;
 wire \mem[29][5] ;
 wire \mem[29][6] ;
 wire \mem[29][7] ;
 wire \mem[29][8] ;
 wire \mem[29][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[30][0] ;
 wire \mem[30][10] ;
 wire \mem[30][11] ;
 wire \mem[30][12] ;
 wire \mem[30][13] ;
 wire \mem[30][14] ;
 wire \mem[30][15] ;
 wire \mem[30][16] ;
 wire \mem[30][17] ;
 wire \mem[30][18] ;
 wire \mem[30][19] ;
 wire \mem[30][1] ;
 wire \mem[30][20] ;
 wire \mem[30][21] ;
 wire \mem[30][22] ;
 wire \mem[30][23] ;
 wire \mem[30][24] ;
 wire \mem[30][25] ;
 wire \mem[30][26] ;
 wire \mem[30][27] ;
 wire \mem[30][28] ;
 wire \mem[30][29] ;
 wire \mem[30][2] ;
 wire \mem[30][30] ;
 wire \mem[30][31] ;
 wire \mem[30][3] ;
 wire \mem[30][4] ;
 wire \mem[30][5] ;
 wire \mem[30][6] ;
 wire \mem[30][7] ;
 wire \mem[30][8] ;
 wire \mem[30][9] ;
 wire \mem[31][0] ;
 wire \mem[31][10] ;
 wire \mem[31][11] ;
 wire \mem[31][12] ;
 wire \mem[31][13] ;
 wire \mem[31][14] ;
 wire \mem[31][15] ;
 wire \mem[31][16] ;
 wire \mem[31][17] ;
 wire \mem[31][18] ;
 wire \mem[31][19] ;
 wire \mem[31][1] ;
 wire \mem[31][20] ;
 wire \mem[31][21] ;
 wire \mem[31][22] ;
 wire \mem[31][23] ;
 wire \mem[31][24] ;
 wire \mem[31][25] ;
 wire \mem[31][26] ;
 wire \mem[31][27] ;
 wire \mem[31][28] ;
 wire \mem[31][29] ;
 wire \mem[31][2] ;
 wire \mem[31][30] ;
 wire \mem[31][31] ;
 wire \mem[31][3] ;
 wire \mem[31][4] ;
 wire \mem[31][5] ;
 wire \mem[31][6] ;
 wire \mem[31][7] ;
 wire \mem[31][8] ;
 wire \mem[31][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;

 sky130_fd_sc_hd__clkbuf_2 _4317_ (.A(net7),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_2 _4318_ (.A(net6),
    .X(_0993_));
 sky130_fd_sc_hd__and2b_1 _4319_ (.A_N(net8),
    .B(net9),
    .X(_0994_));
 sky130_fd_sc_hd__buf_2 _4320_ (.A(net10),
    .X(_0995_));
 sky130_fd_sc_hd__and4b_2 _4321_ (.A_N(_0992_),
    .B(_0993_),
    .C(_0994_),
    .D(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__buf_4 _4322_ (.A(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__buf_2 _4323_ (.A(net9),
    .X(_0998_));
 sky130_fd_sc_hd__buf_2 _4324_ (.A(net8),
    .X(_0999_));
 sky130_fd_sc_hd__and2_2 _4325_ (.A(_0998_),
    .B(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__clkbuf_4 _4326_ (.A(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__nor3_1 _4327_ (.A(net10),
    .B(net7),
    .C(net6),
    .Y(_1002_));
 sky130_fd_sc_hd__clkbuf_4 _4328_ (.A(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__buf_4 _4329_ (.A(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__and3_1 _4330_ (.A(\mem[12][19] ),
    .B(_1001_),
    .C(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__buf_4 _4331_ (.A(_0995_),
    .X(_1006_));
 sky130_fd_sc_hd__and4b_4 _4332_ (.A_N(net7),
    .B(net6),
    .C(_0998_),
    .D(_0999_),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_4 _4333_ (.A(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__and3_1 _4334_ (.A(\mem[29][19] ),
    .B(_1006_),
    .C(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__buf_2 _4335_ (.A(net10),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_4 _4336_ (.A(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__and4b_2 _4337_ (.A_N(_0993_),
    .B(_0998_),
    .C(_0999_),
    .D(net7),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_4 _4338_ (.A(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__and3_1 _4339_ (.A(\mem[30][19] ),
    .B(_1011_),
    .C(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__a2111o_1 _4340_ (.A1(\mem[25][19] ),
    .A2(_0997_),
    .B1(_1005_),
    .C1(_1009_),
    .D1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and4bb_2 _4341_ (.A_N(_0995_),
    .B_N(_0993_),
    .C(_0994_),
    .D(_0992_),
    .X(_1016_));
 sky130_fd_sc_hd__buf_4 _4342_ (.A(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__clkinv_2 _4343_ (.A(net10),
    .Y(_1018_));
 sky130_fd_sc_hd__clkbuf_4 _4344_ (.A(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__and3_1 _4345_ (.A(\mem[13][19] ),
    .B(_1019_),
    .C(_1007_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_4 _4346_ (.A(_0994_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_4 _4347_ (.A(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__nor3b_1 _4348_ (.A(net7),
    .B(net6),
    .C_N(net10),
    .Y(_1023_));
 sky130_fd_sc_hd__clkbuf_4 _4349_ (.A(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__and3_1 _4350_ (.A(\mem[24][19] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__buf_4 _4351_ (.A(_1018_),
    .X(_1026_));
 sky130_fd_sc_hd__and4_4 _4352_ (.A(_0992_),
    .B(net6),
    .C(_0998_),
    .D(_0999_),
    .X(_1027_));
 sky130_fd_sc_hd__buf_4 _4353_ (.A(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__and3_1 _4354_ (.A(\mem[15][19] ),
    .B(_1026_),
    .C(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__a2111o_1 _4355_ (.A1(\mem[10][19] ),
    .A2(_1017_),
    .B1(_1020_),
    .C1(_1025_),
    .D1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__inv_2 _4356_ (.A(\mem[3][19] ),
    .Y(_1031_));
 sky130_fd_sc_hd__or4bb_4 _4357_ (.A(net9),
    .B(net8),
    .C_N(net7),
    .D_N(net6),
    .X(_1032_));
 sky130_fd_sc_hd__or2_1 _4358_ (.A(_0995_),
    .B(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4359_ (.A(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_4 _4360_ (.A(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_4 _4361_ (.A(_1010_),
    .X(_1036_));
 sky130_fd_sc_hd__or4b_4 _4362_ (.A(net7),
    .B(_0998_),
    .C(_0999_),
    .D_N(net6),
    .X(_1037_));
 sky130_fd_sc_hd__or3b_1 _4363_ (.A(_1036_),
    .B(_1037_),
    .C_N(\mem[1][19] ),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_4 _4364_ (.A(_1010_),
    .X(_1039_));
 sky130_fd_sc_hd__or4bb_4 _4365_ (.A(net7),
    .B(_0998_),
    .C_N(_0999_),
    .D_N(net6),
    .X(_1040_));
 sky130_fd_sc_hd__clkbuf_4 _4366_ (.A(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__or3b_1 _4367_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][19] ),
    .X(_1042_));
 sky130_fd_sc_hd__inv_2 _4368_ (.A(\mem[19][19] ),
    .Y(_1043_));
 sky130_fd_sc_hd__buf_2 _4369_ (.A(_1018_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_4 _4370_ (.A(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__clkbuf_4 _4371_ (.A(_1032_),
    .X(_1046_));
 sky130_fd_sc_hd__or3_1 _4372_ (.A(_1043_),
    .B(_1045_),
    .C(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__o2111ai_1 _4373_ (.A1(_1031_),
    .A2(_1035_),
    .B1(_1038_),
    .C1(_1042_),
    .D1(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__or4b_1 _4374_ (.A(net6),
    .B(_0998_),
    .C(_0999_),
    .D_N(net7),
    .X(_1049_));
 sky130_fd_sc_hd__nor2_2 _4375_ (.A(_1044_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__buf_4 _4376_ (.A(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_4 _4377_ (.A(_1003_),
    .X(_1052_));
 sky130_fd_sc_hd__and2b_1 _4378_ (.A_N(_0998_),
    .B(_0999_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_4 _4379_ (.A(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_4 _4380_ (.A(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__and3_1 _4381_ (.A(\mem[4][19] ),
    .B(_1052_),
    .C(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_4 _4382_ (.A(_1010_),
    .X(_1057_));
 sky130_fd_sc_hd__and4bb_4 _4383_ (.A_N(_0993_),
    .B_N(_0998_),
    .C(_0999_),
    .D(_0992_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_4 _4384_ (.A(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__and3_1 _4385_ (.A(\mem[22][19] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_4 _4386_ (.A(_1054_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_4 _4387_ (.A(_1023_),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_4 _4388_ (.A(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__and3_1 _4389_ (.A(\mem[20][19] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__a2111o_1 _4390_ (.A1(\mem[18][19] ),
    .A2(_1051_),
    .B1(_1056_),
    .C1(_1060_),
    .D1(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__or4_1 _4391_ (.A(_1015_),
    .B(_1030_),
    .C(_1048_),
    .D(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_4 _4392_ (.A(net10),
    .X(_1067_));
 sky130_fd_sc_hd__and4b_2 _4393_ (.A_N(_0993_),
    .B(_1021_),
    .C(_1067_),
    .D(_0992_),
    .X(_1068_));
 sky130_fd_sc_hd__buf_4 _4394_ (.A(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__and4_4 _4395_ (.A(_1010_),
    .B(_0992_),
    .C(_0993_),
    .D(_1021_),
    .X(_1070_));
 sky130_fd_sc_hd__and2_2 _4396_ (.A(_1000_),
    .B(_1062_),
    .X(_1071_));
 sky130_fd_sc_hd__a22o_1 _4397_ (.A1(\mem[27][19] ),
    .A2(_1070_),
    .B1(_1071_),
    .B2(\mem[28][19] ),
    .X(_1072_));
 sky130_fd_sc_hd__buf_4 _4398_ (.A(_1067_),
    .X(_1073_));
 sky130_fd_sc_hd__and2_2 _4399_ (.A(_1044_),
    .B(_1012_),
    .X(_1074_));
 sky130_fd_sc_hd__a32o_1 _4400_ (.A1(_1073_),
    .A2(\mem[31][19] ),
    .A3(_1028_),
    .B1(_1074_),
    .B2(\mem[14][19] ),
    .X(_1075_));
 sky130_fd_sc_hd__and4bb_4 _4401_ (.A_N(_1010_),
    .B_N(_0992_),
    .C(_0993_),
    .D(_1021_),
    .X(_1076_));
 sky130_fd_sc_hd__buf_4 _4402_ (.A(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__and4_2 _4403_ (.A(_1044_),
    .B(_0992_),
    .C(_0993_),
    .D(_1021_),
    .X(_1078_));
 sky130_fd_sc_hd__buf_4 _4404_ (.A(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__a22o_1 _4405_ (.A1(\mem[9][19] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][19] ),
    .X(_1080_));
 sky130_fd_sc_hd__a2111o_1 _4406_ (.A1(\mem[26][19] ),
    .A2(_1069_),
    .B1(_1072_),
    .C1(_1075_),
    .D1(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__and2_2 _4407_ (.A(_1022_),
    .B(_1052_),
    .X(_1082_));
 sky130_fd_sc_hd__buf_4 _4408_ (.A(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__and2_1 _4409_ (.A(_1045_),
    .B(_1059_),
    .X(_1084_));
 sky130_fd_sc_hd__buf_4 _4410_ (.A(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__nor3b_4 _4411_ (.A(_0998_),
    .B(_0999_),
    .C_N(_1062_),
    .Y(_1086_));
 sky130_fd_sc_hd__buf_4 _4412_ (.A(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__and4_2 _4413_ (.A(_1044_),
    .B(_0992_),
    .C(_0993_),
    .D(_1054_),
    .X(_1088_));
 sky130_fd_sc_hd__buf_4 _4414_ (.A(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__a22o_1 _4415_ (.A1(\mem[16][19] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][19] ),
    .X(_1090_));
 sky130_fd_sc_hd__a221o_1 _4416_ (.A1(\mem[8][19] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][19] ),
    .C1(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__nor2_2 _4417_ (.A(_1011_),
    .B(_1049_),
    .Y(_1092_));
 sky130_fd_sc_hd__buf_4 _4418_ (.A(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__and4_2 _4419_ (.A(_1073_),
    .B(_0992_),
    .C(_0993_),
    .D(_1061_),
    .X(_1094_));
 sky130_fd_sc_hd__buf_4 _4420_ (.A(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__nor2_2 _4421_ (.A(_1026_),
    .B(_1040_),
    .Y(_1096_));
 sky130_fd_sc_hd__buf_4 _4422_ (.A(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_2 _4423_ (.A(_1026_),
    .B(_1037_),
    .Y(_1098_));
 sky130_fd_sc_hd__buf_4 _4424_ (.A(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_1 _4425_ (.A1(\mem[21][19] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][19] ),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _4426_ (.A1(\mem[2][19] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][19] ),
    .C1(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__or4_4 _4427_ (.A(_1066_),
    .B(_1081_),
    .C(_1091_),
    .D(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _4428_ (.A(_1102_),
    .X(net92));
 sky130_fd_sc_hd__and3_1 _4429_ (.A(\mem[12][20] ),
    .B(_1001_),
    .C(_1004_),
    .X(_1103_));
 sky130_fd_sc_hd__and3_1 _4430_ (.A(\mem[29][20] ),
    .B(_1006_),
    .C(_1008_),
    .X(_1104_));
 sky130_fd_sc_hd__and3_1 _4431_ (.A(\mem[30][20] ),
    .B(_1011_),
    .C(_1013_),
    .X(_1105_));
 sky130_fd_sc_hd__a2111o_1 _4432_ (.A1(\mem[25][20] ),
    .A2(_0997_),
    .B1(_1103_),
    .C1(_1104_),
    .D1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__buf_2 _4433_ (.A(_1018_),
    .X(_1107_));
 sky130_fd_sc_hd__and3_1 _4434_ (.A(\mem[15][20] ),
    .B(_1107_),
    .C(_1028_),
    .X(_1108_));
 sky130_fd_sc_hd__and3_1 _4435_ (.A(\mem[24][20] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1109_));
 sky130_fd_sc_hd__buf_2 _4436_ (.A(_1007_),
    .X(_1110_));
 sky130_fd_sc_hd__and3_1 _4437_ (.A(\mem[13][20] ),
    .B(_1026_),
    .C(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__a2111o_1 _4438_ (.A1(\mem[10][20] ),
    .A2(_1017_),
    .B1(_1108_),
    .C1(_1109_),
    .D1(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(\mem[3][20] ),
    .Y(_1113_));
 sky130_fd_sc_hd__inv_2 _4440_ (.A(\mem[19][20] ),
    .Y(_1114_));
 sky130_fd_sc_hd__clkbuf_4 _4441_ (.A(_1044_),
    .X(_1115_));
 sky130_fd_sc_hd__or3_1 _4442_ (.A(_1114_),
    .B(_1115_),
    .C(_1046_),
    .X(_1116_));
 sky130_fd_sc_hd__or3b_1 _4443_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][20] ),
    .X(_1117_));
 sky130_fd_sc_hd__buf_2 _4444_ (.A(_1010_),
    .X(_1118_));
 sky130_fd_sc_hd__buf_2 _4445_ (.A(_1037_),
    .X(_1119_));
 sky130_fd_sc_hd__or3b_1 _4446_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][20] ),
    .X(_1120_));
 sky130_fd_sc_hd__o2111ai_1 _4447_ (.A1(_1113_),
    .A2(_1035_),
    .B1(_1116_),
    .C1(_1117_),
    .D1(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__and3_1 _4448_ (.A(\mem[4][20] ),
    .B(_1052_),
    .C(_1055_),
    .X(_1122_));
 sky130_fd_sc_hd__and3_1 _4449_ (.A(\mem[22][20] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1123_));
 sky130_fd_sc_hd__and3_1 _4450_ (.A(\mem[20][20] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1124_));
 sky130_fd_sc_hd__a2111o_1 _4451_ (.A1(\mem[18][20] ),
    .A2(_1051_),
    .B1(_1122_),
    .C1(_1123_),
    .D1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__or4_1 _4452_ (.A(_1106_),
    .B(_1112_),
    .C(_1121_),
    .D(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__a22o_1 _4453_ (.A1(\mem[9][20] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][20] ),
    .X(_1127_));
 sky130_fd_sc_hd__buf_4 _4454_ (.A(_1070_),
    .X(_1128_));
 sky130_fd_sc_hd__buf_4 _4455_ (.A(_1071_),
    .X(_1129_));
 sky130_fd_sc_hd__a22o_1 _4456_ (.A1(\mem[27][20] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][20] ),
    .X(_1130_));
 sky130_fd_sc_hd__buf_4 _4457_ (.A(_1073_),
    .X(_1131_));
 sky130_fd_sc_hd__buf_4 _4458_ (.A(_1028_),
    .X(_1132_));
 sky130_fd_sc_hd__buf_4 _4459_ (.A(_1074_),
    .X(_1133_));
 sky130_fd_sc_hd__a32o_1 _4460_ (.A1(\mem[31][20] ),
    .A2(_1131_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][20] ),
    .X(_1134_));
 sky130_fd_sc_hd__a2111o_1 _4461_ (.A1(\mem[26][20] ),
    .A2(_1069_),
    .B1(_1127_),
    .C1(_1130_),
    .D1(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__a22o_1 _4462_ (.A1(\mem[16][20] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][20] ),
    .X(_1136_));
 sky130_fd_sc_hd__a221o_1 _4463_ (.A1(\mem[8][20] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][20] ),
    .C1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__a22o_1 _4464_ (.A1(\mem[21][20] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][20] ),
    .X(_1138_));
 sky130_fd_sc_hd__a221o_1 _4465_ (.A1(\mem[2][20] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][20] ),
    .C1(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__or4_4 _4466_ (.A(_1126_),
    .B(_1135_),
    .C(_1137_),
    .D(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _4467_ (.A(_1140_),
    .X(net94));
 sky130_fd_sc_hd__and3_1 _4468_ (.A(\mem[12][21] ),
    .B(_1001_),
    .C(_1004_),
    .X(_1141_));
 sky130_fd_sc_hd__and3_1 _4469_ (.A(\mem[29][21] ),
    .B(_1006_),
    .C(_1008_),
    .X(_1142_));
 sky130_fd_sc_hd__and3_1 _4470_ (.A(\mem[30][21] ),
    .B(_1011_),
    .C(_1013_),
    .X(_1143_));
 sky130_fd_sc_hd__a2111o_1 _4471_ (.A1(\mem[25][21] ),
    .A2(_0997_),
    .B1(_1141_),
    .C1(_1142_),
    .D1(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__and3_1 _4472_ (.A(\mem[15][21] ),
    .B(_1107_),
    .C(_1028_),
    .X(_1145_));
 sky130_fd_sc_hd__and3_1 _4473_ (.A(\mem[24][21] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1146_));
 sky130_fd_sc_hd__buf_2 _4474_ (.A(_1044_),
    .X(_1147_));
 sky130_fd_sc_hd__and3_1 _4475_ (.A(\mem[13][21] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1148_));
 sky130_fd_sc_hd__a2111o_1 _4476_ (.A1(\mem[10][21] ),
    .A2(_1017_),
    .B1(_1145_),
    .C1(_1146_),
    .D1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__inv_2 _4477_ (.A(\mem[3][21] ),
    .Y(_1150_));
 sky130_fd_sc_hd__inv_2 _4478_ (.A(\mem[19][21] ),
    .Y(_1151_));
 sky130_fd_sc_hd__clkbuf_4 _4479_ (.A(_1032_),
    .X(_1152_));
 sky130_fd_sc_hd__or3_1 _4480_ (.A(_1151_),
    .B(_1115_),
    .C(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__or3b_1 _4481_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][21] ),
    .X(_1154_));
 sky130_fd_sc_hd__or3b_1 _4482_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][21] ),
    .X(_1155_));
 sky130_fd_sc_hd__o2111ai_1 _4483_ (.A1(_1150_),
    .A2(_1035_),
    .B1(_1153_),
    .C1(_1154_),
    .D1(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__and3_1 _4484_ (.A(\mem[4][21] ),
    .B(_1052_),
    .C(_1055_),
    .X(_1157_));
 sky130_fd_sc_hd__and3_1 _4485_ (.A(\mem[22][21] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1158_));
 sky130_fd_sc_hd__and3_1 _4486_ (.A(\mem[20][21] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1159_));
 sky130_fd_sc_hd__a2111o_1 _4487_ (.A1(\mem[18][21] ),
    .A2(_1051_),
    .B1(_1157_),
    .C1(_1158_),
    .D1(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__or4_1 _4488_ (.A(_1144_),
    .B(_1149_),
    .C(_1156_),
    .D(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__a22o_1 _4489_ (.A1(\mem[9][21] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][21] ),
    .X(_1162_));
 sky130_fd_sc_hd__a22o_1 _4490_ (.A1(\mem[27][21] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][21] ),
    .X(_1163_));
 sky130_fd_sc_hd__a32o_1 _4491_ (.A1(\mem[31][21] ),
    .A2(_1131_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][21] ),
    .X(_1164_));
 sky130_fd_sc_hd__a2111o_1 _4492_ (.A1(\mem[26][21] ),
    .A2(_1069_),
    .B1(_1162_),
    .C1(_1163_),
    .D1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__a22o_1 _4493_ (.A1(\mem[16][21] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][21] ),
    .X(_1166_));
 sky130_fd_sc_hd__a221o_1 _4494_ (.A1(\mem[8][21] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][21] ),
    .C1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__a22o_1 _4495_ (.A1(\mem[21][21] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][21] ),
    .X(_1168_));
 sky130_fd_sc_hd__a221o_1 _4496_ (.A1(\mem[2][21] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][21] ),
    .C1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__or4_4 _4497_ (.A(_1161_),
    .B(_1165_),
    .C(_1167_),
    .D(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__clkbuf_1 _4498_ (.A(_1170_),
    .X(net95));
 sky130_fd_sc_hd__and3_1 _4499_ (.A(\mem[12][22] ),
    .B(_1001_),
    .C(_1004_),
    .X(_1171_));
 sky130_fd_sc_hd__and3_1 _4500_ (.A(\mem[29][22] ),
    .B(_1006_),
    .C(_1008_),
    .X(_1172_));
 sky130_fd_sc_hd__and3_1 _4501_ (.A(\mem[30][22] ),
    .B(_1011_),
    .C(_1013_),
    .X(_1173_));
 sky130_fd_sc_hd__a2111o_1 _4502_ (.A1(\mem[25][22] ),
    .A2(_0997_),
    .B1(_1171_),
    .C1(_1172_),
    .D1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__and3_1 _4503_ (.A(\mem[15][22] ),
    .B(_1107_),
    .C(_1028_),
    .X(_1175_));
 sky130_fd_sc_hd__and3_1 _4504_ (.A(\mem[24][22] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1176_));
 sky130_fd_sc_hd__and3_1 _4505_ (.A(\mem[13][22] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1177_));
 sky130_fd_sc_hd__a2111o_1 _4506_ (.A1(\mem[10][22] ),
    .A2(_1017_),
    .B1(_1175_),
    .C1(_1176_),
    .D1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__inv_2 _4507_ (.A(\mem[3][22] ),
    .Y(_1179_));
 sky130_fd_sc_hd__clkbuf_4 _4508_ (.A(_1040_),
    .X(_1180_));
 sky130_fd_sc_hd__or3b_1 _4509_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][22] ),
    .X(_1181_));
 sky130_fd_sc_hd__inv_2 _4510_ (.A(\mem[19][22] ),
    .Y(_1182_));
 sky130_fd_sc_hd__or3_1 _4511_ (.A(_1182_),
    .B(_1045_),
    .C(_1046_),
    .X(_1183_));
 sky130_fd_sc_hd__or3b_1 _4512_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][22] ),
    .X(_1184_));
 sky130_fd_sc_hd__o2111ai_2 _4513_ (.A1(_1179_),
    .A2(_1035_),
    .B1(_1181_),
    .C1(_1183_),
    .D1(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__and3_1 _4514_ (.A(\mem[4][22] ),
    .B(_1052_),
    .C(_1055_),
    .X(_1186_));
 sky130_fd_sc_hd__and3_1 _4515_ (.A(\mem[22][22] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1187_));
 sky130_fd_sc_hd__and3_1 _4516_ (.A(\mem[20][22] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1188_));
 sky130_fd_sc_hd__a2111o_1 _4517_ (.A1(\mem[18][22] ),
    .A2(_1051_),
    .B1(_1186_),
    .C1(_1187_),
    .D1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__or4_1 _4518_ (.A(_1174_),
    .B(_1178_),
    .C(_1185_),
    .D(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__a22o_1 _4519_ (.A1(\mem[9][22] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][22] ),
    .X(_1191_));
 sky130_fd_sc_hd__a22o_1 _4520_ (.A1(\mem[27][22] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][22] ),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_4 _4521_ (.A(_1073_),
    .X(_1193_));
 sky130_fd_sc_hd__a32o_1 _4522_ (.A1(\mem[31][22] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][22] ),
    .X(_1194_));
 sky130_fd_sc_hd__a2111o_1 _4523_ (.A1(\mem[26][22] ),
    .A2(_1069_),
    .B1(_1191_),
    .C1(_1192_),
    .D1(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_1 _4524_ (.A1(\mem[16][22] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][22] ),
    .X(_1196_));
 sky130_fd_sc_hd__a221o_1 _4525_ (.A1(\mem[8][22] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][22] ),
    .C1(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__a22o_1 _4526_ (.A1(\mem[21][22] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][22] ),
    .X(_1198_));
 sky130_fd_sc_hd__a221o_1 _4527_ (.A1(\mem[2][22] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][22] ),
    .C1(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__or4_4 _4528_ (.A(_1190_),
    .B(_1195_),
    .C(_1197_),
    .D(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _4529_ (.A(_1200_),
    .X(net96));
 sky130_fd_sc_hd__and3_1 _4530_ (.A(\mem[12][23] ),
    .B(_1001_),
    .C(_1004_),
    .X(_1201_));
 sky130_fd_sc_hd__buf_4 _4531_ (.A(_0995_),
    .X(_1202_));
 sky130_fd_sc_hd__and3_1 _4532_ (.A(\mem[29][23] ),
    .B(_1202_),
    .C(_1008_),
    .X(_1203_));
 sky130_fd_sc_hd__and3_1 _4533_ (.A(\mem[30][23] ),
    .B(_1011_),
    .C(_1013_),
    .X(_1204_));
 sky130_fd_sc_hd__a2111o_1 _4534_ (.A1(\mem[25][23] ),
    .A2(_0997_),
    .B1(_1201_),
    .C1(_1203_),
    .D1(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__and3_1 _4535_ (.A(\mem[15][23] ),
    .B(_1107_),
    .C(_1028_),
    .X(_1206_));
 sky130_fd_sc_hd__and3_1 _4536_ (.A(\mem[24][23] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1207_));
 sky130_fd_sc_hd__and3_1 _4537_ (.A(\mem[13][23] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1208_));
 sky130_fd_sc_hd__a2111o_1 _4538_ (.A1(\mem[10][23] ),
    .A2(_1017_),
    .B1(_1206_),
    .C1(_1207_),
    .D1(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__inv_2 _4539_ (.A(\mem[3][23] ),
    .Y(_1210_));
 sky130_fd_sc_hd__inv_2 _4540_ (.A(\mem[19][23] ),
    .Y(_1211_));
 sky130_fd_sc_hd__or3_1 _4541_ (.A(_1211_),
    .B(_1115_),
    .C(_1152_),
    .X(_1212_));
 sky130_fd_sc_hd__or3b_1 _4542_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][23] ),
    .X(_1213_));
 sky130_fd_sc_hd__or3b_1 _4543_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][23] ),
    .X(_1214_));
 sky130_fd_sc_hd__o2111ai_1 _4544_ (.A1(_1210_),
    .A2(_1035_),
    .B1(_1212_),
    .C1(_1213_),
    .D1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__and3_1 _4545_ (.A(\mem[4][23] ),
    .B(_1052_),
    .C(_1055_),
    .X(_1216_));
 sky130_fd_sc_hd__and3_1 _4546_ (.A(\mem[22][23] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1217_));
 sky130_fd_sc_hd__and3_1 _4547_ (.A(\mem[20][23] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1218_));
 sky130_fd_sc_hd__a2111o_1 _4548_ (.A1(\mem[18][23] ),
    .A2(_1051_),
    .B1(_1216_),
    .C1(_1217_),
    .D1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__or4_1 _4549_ (.A(_1205_),
    .B(_1209_),
    .C(_1215_),
    .D(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__a22o_1 _4550_ (.A1(\mem[9][23] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][23] ),
    .X(_1221_));
 sky130_fd_sc_hd__a22o_1 _4551_ (.A1(\mem[27][23] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][23] ),
    .X(_1222_));
 sky130_fd_sc_hd__a32o_1 _4552_ (.A1(\mem[31][23] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][23] ),
    .X(_1223_));
 sky130_fd_sc_hd__a2111o_1 _4553_ (.A1(\mem[26][23] ),
    .A2(_1069_),
    .B1(_1221_),
    .C1(_1222_),
    .D1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a22o_1 _4554_ (.A1(\mem[16][23] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][23] ),
    .X(_1225_));
 sky130_fd_sc_hd__a221o_1 _4555_ (.A1(\mem[8][23] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][23] ),
    .C1(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__a22o_1 _4556_ (.A1(\mem[21][23] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][23] ),
    .X(_1227_));
 sky130_fd_sc_hd__a221o_1 _4557_ (.A1(\mem[2][23] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][23] ),
    .C1(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__or4_4 _4558_ (.A(_1220_),
    .B(_1224_),
    .C(_1226_),
    .D(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _4559_ (.A(_1229_),
    .X(net97));
 sky130_fd_sc_hd__and3_1 _4560_ (.A(\mem[12][24] ),
    .B(_1001_),
    .C(_1004_),
    .X(_1230_));
 sky130_fd_sc_hd__and3_1 _4561_ (.A(\mem[29][24] ),
    .B(_1202_),
    .C(_1008_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_4 _4562_ (.A(_0995_),
    .X(_1232_));
 sky130_fd_sc_hd__and3_1 _4563_ (.A(\mem[30][24] ),
    .B(_1232_),
    .C(_1013_),
    .X(_1233_));
 sky130_fd_sc_hd__a2111o_1 _4564_ (.A1(\mem[25][24] ),
    .A2(_0997_),
    .B1(_1230_),
    .C1(_1231_),
    .D1(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__buf_4 _4565_ (.A(_1027_),
    .X(_1235_));
 sky130_fd_sc_hd__and3_1 _4566_ (.A(\mem[15][24] ),
    .B(_1107_),
    .C(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__and3_1 _4567_ (.A(\mem[24][24] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1237_));
 sky130_fd_sc_hd__and3_1 _4568_ (.A(\mem[13][24] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1238_));
 sky130_fd_sc_hd__a2111o_1 _4569_ (.A1(\mem[10][24] ),
    .A2(_1017_),
    .B1(_1236_),
    .C1(_1237_),
    .D1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__inv_2 _4570_ (.A(\mem[3][24] ),
    .Y(_1240_));
 sky130_fd_sc_hd__or3b_1 _4571_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][24] ),
    .X(_1241_));
 sky130_fd_sc_hd__inv_2 _4572_ (.A(\mem[19][24] ),
    .Y(_1242_));
 sky130_fd_sc_hd__or3_1 _4573_ (.A(_1242_),
    .B(_1045_),
    .C(_1046_),
    .X(_1243_));
 sky130_fd_sc_hd__or3b_1 _4574_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][24] ),
    .X(_1244_));
 sky130_fd_sc_hd__o2111ai_1 _4575_ (.A1(_1240_),
    .A2(_1035_),
    .B1(_1241_),
    .C1(_1243_),
    .D1(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__and3_1 _4576_ (.A(\mem[4][24] ),
    .B(_1052_),
    .C(_1055_),
    .X(_1246_));
 sky130_fd_sc_hd__and3_1 _4577_ (.A(\mem[22][24] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1247_));
 sky130_fd_sc_hd__and3_1 _4578_ (.A(\mem[20][24] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1248_));
 sky130_fd_sc_hd__a2111o_1 _4579_ (.A1(\mem[18][24] ),
    .A2(_1051_),
    .B1(_1246_),
    .C1(_1247_),
    .D1(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__or4_1 _4580_ (.A(_1234_),
    .B(_1239_),
    .C(_1245_),
    .D(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__a22o_1 _4581_ (.A1(\mem[9][24] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][24] ),
    .X(_1251_));
 sky130_fd_sc_hd__a22o_1 _4582_ (.A1(\mem[27][24] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][24] ),
    .X(_1252_));
 sky130_fd_sc_hd__a32o_1 _4583_ (.A1(\mem[31][24] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][24] ),
    .X(_1253_));
 sky130_fd_sc_hd__a2111o_1 _4584_ (.A1(\mem[26][24] ),
    .A2(_1069_),
    .B1(_1251_),
    .C1(_1252_),
    .D1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a22o_1 _4585_ (.A1(\mem[16][24] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][24] ),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_1 _4586_ (.A1(\mem[8][24] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][24] ),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__a22o_1 _4587_ (.A1(\mem[21][24] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][24] ),
    .X(_1257_));
 sky130_fd_sc_hd__a221o_1 _4588_ (.A1(\mem[2][24] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][24] ),
    .C1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__or4_1 _4589_ (.A(_1250_),
    .B(_1254_),
    .C(_1256_),
    .D(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__buf_6 _4590_ (.A(_1259_),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 _4591_ (.A(_1003_),
    .X(_1260_));
 sky130_fd_sc_hd__and3_1 _4592_ (.A(\mem[12][25] ),
    .B(_1001_),
    .C(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__and3_1 _4593_ (.A(\mem[29][25] ),
    .B(_1202_),
    .C(_1008_),
    .X(_1262_));
 sky130_fd_sc_hd__and3_1 _4594_ (.A(\mem[30][25] ),
    .B(_1232_),
    .C(_1013_),
    .X(_1263_));
 sky130_fd_sc_hd__a2111o_1 _4595_ (.A1(\mem[25][25] ),
    .A2(_0997_),
    .B1(_1261_),
    .C1(_1262_),
    .D1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__and3_1 _4596_ (.A(\mem[15][25] ),
    .B(_1107_),
    .C(_1235_),
    .X(_1265_));
 sky130_fd_sc_hd__and3_1 _4597_ (.A(\mem[24][25] ),
    .B(_1022_),
    .C(_1024_),
    .X(_1266_));
 sky130_fd_sc_hd__and3_1 _4598_ (.A(\mem[13][25] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1267_));
 sky130_fd_sc_hd__a2111o_1 _4599_ (.A1(\mem[10][25] ),
    .A2(_1017_),
    .B1(_1265_),
    .C1(_1266_),
    .D1(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__inv_2 _4600_ (.A(\mem[3][25] ),
    .Y(_1269_));
 sky130_fd_sc_hd__or3b_1 _4601_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][25] ),
    .X(_1270_));
 sky130_fd_sc_hd__inv_2 _4602_ (.A(\mem[19][25] ),
    .Y(_1271_));
 sky130_fd_sc_hd__or3_1 _4603_ (.A(_1271_),
    .B(_1045_),
    .C(_1046_),
    .X(_1272_));
 sky130_fd_sc_hd__or3b_1 _4604_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][25] ),
    .X(_1273_));
 sky130_fd_sc_hd__o2111ai_1 _4605_ (.A1(_1269_),
    .A2(_1035_),
    .B1(_1270_),
    .C1(_1272_),
    .D1(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__buf_4 _4606_ (.A(_1053_),
    .X(_1275_));
 sky130_fd_sc_hd__and3_1 _4607_ (.A(\mem[4][25] ),
    .B(_1052_),
    .C(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__and3_1 _4608_ (.A(\mem[22][25] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1277_));
 sky130_fd_sc_hd__and3_1 _4609_ (.A(\mem[20][25] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1278_));
 sky130_fd_sc_hd__a2111o_1 _4610_ (.A1(\mem[18][25] ),
    .A2(_1051_),
    .B1(_1276_),
    .C1(_1277_),
    .D1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__or4_1 _4611_ (.A(_1264_),
    .B(_1268_),
    .C(_1274_),
    .D(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__a22o_1 _4612_ (.A1(\mem[9][25] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][25] ),
    .X(_1281_));
 sky130_fd_sc_hd__a22o_1 _4613_ (.A1(\mem[27][25] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][25] ),
    .X(_1282_));
 sky130_fd_sc_hd__a32o_1 _4614_ (.A1(\mem[31][25] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][25] ),
    .X(_1283_));
 sky130_fd_sc_hd__a2111o_1 _4615_ (.A1(\mem[26][25] ),
    .A2(_1069_),
    .B1(_1281_),
    .C1(_1282_),
    .D1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a22o_1 _4616_ (.A1(\mem[16][25] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][25] ),
    .X(_1285_));
 sky130_fd_sc_hd__a221o_1 _4617_ (.A1(\mem[8][25] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][25] ),
    .C1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__a22o_1 _4618_ (.A1(\mem[21][25] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][25] ),
    .X(_1287_));
 sky130_fd_sc_hd__a221o_1 _4619_ (.A1(\mem[2][25] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][25] ),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__or4_4 _4620_ (.A(_1280_),
    .B(_1284_),
    .C(_1286_),
    .D(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _4621_ (.A(_1289_),
    .X(net99));
 sky130_fd_sc_hd__and3_1 _4622_ (.A(\mem[12][26] ),
    .B(_1001_),
    .C(_1260_),
    .X(_1290_));
 sky130_fd_sc_hd__and3_1 _4623_ (.A(\mem[29][26] ),
    .B(_1202_),
    .C(_1008_),
    .X(_1291_));
 sky130_fd_sc_hd__and3_1 _4624_ (.A(\mem[30][26] ),
    .B(_1232_),
    .C(_1013_),
    .X(_1292_));
 sky130_fd_sc_hd__a2111o_1 _4625_ (.A1(\mem[25][26] ),
    .A2(_0997_),
    .B1(_1290_),
    .C1(_1291_),
    .D1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__and3_1 _4626_ (.A(\mem[15][26] ),
    .B(_1107_),
    .C(_1235_),
    .X(_1294_));
 sky130_fd_sc_hd__buf_4 _4627_ (.A(_1023_),
    .X(_1295_));
 sky130_fd_sc_hd__and3_1 _4628_ (.A(\mem[24][26] ),
    .B(_1022_),
    .C(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__and3_1 _4629_ (.A(\mem[13][26] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1297_));
 sky130_fd_sc_hd__a2111o_1 _4630_ (.A1(\mem[10][26] ),
    .A2(_1017_),
    .B1(_1294_),
    .C1(_1296_),
    .D1(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__inv_2 _4631_ (.A(\mem[3][26] ),
    .Y(_1299_));
 sky130_fd_sc_hd__inv_2 _4632_ (.A(\mem[19][26] ),
    .Y(_1300_));
 sky130_fd_sc_hd__or3_1 _4633_ (.A(_1300_),
    .B(_1115_),
    .C(_1152_),
    .X(_1301_));
 sky130_fd_sc_hd__or3b_1 _4634_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][26] ),
    .X(_1302_));
 sky130_fd_sc_hd__or3b_1 _4635_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][26] ),
    .X(_1303_));
 sky130_fd_sc_hd__o2111ai_1 _4636_ (.A1(_1299_),
    .A2(_1035_),
    .B1(_1301_),
    .C1(_1302_),
    .D1(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__and3_1 _4637_ (.A(\mem[4][26] ),
    .B(_1052_),
    .C(_1275_),
    .X(_1305_));
 sky130_fd_sc_hd__and3_1 _4638_ (.A(\mem[22][26] ),
    .B(_1057_),
    .C(_1059_),
    .X(_1306_));
 sky130_fd_sc_hd__and3_1 _4639_ (.A(\mem[20][26] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1307_));
 sky130_fd_sc_hd__a2111o_1 _4640_ (.A1(\mem[18][26] ),
    .A2(_1051_),
    .B1(_1305_),
    .C1(_1306_),
    .D1(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__or4_1 _4641_ (.A(_1293_),
    .B(_1298_),
    .C(_1304_),
    .D(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__a22o_1 _4642_ (.A1(\mem[9][26] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][26] ),
    .X(_1310_));
 sky130_fd_sc_hd__a22o_1 _4643_ (.A1(\mem[27][26] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][26] ),
    .X(_1311_));
 sky130_fd_sc_hd__a32o_1 _4644_ (.A1(\mem[31][26] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][26] ),
    .X(_1312_));
 sky130_fd_sc_hd__a2111o_1 _4645_ (.A1(\mem[26][26] ),
    .A2(_1069_),
    .B1(_1310_),
    .C1(_1311_),
    .D1(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__a22o_1 _4646_ (.A1(\mem[16][26] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][26] ),
    .X(_1314_));
 sky130_fd_sc_hd__a221o_1 _4647_ (.A1(\mem[8][26] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][26] ),
    .C1(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__a22o_1 _4648_ (.A1(\mem[21][26] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][26] ),
    .X(_1316_));
 sky130_fd_sc_hd__a221o_1 _4649_ (.A1(\mem[2][26] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][26] ),
    .C1(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__or4_4 _4650_ (.A(_1309_),
    .B(_1313_),
    .C(_1315_),
    .D(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _4651_ (.A(_1318_),
    .X(net100));
 sky130_fd_sc_hd__buf_4 _4652_ (.A(_1000_),
    .X(_1319_));
 sky130_fd_sc_hd__and3_1 _4653_ (.A(\mem[12][27] ),
    .B(_1319_),
    .C(_1260_),
    .X(_1320_));
 sky130_fd_sc_hd__buf_4 _4654_ (.A(_1007_),
    .X(_1321_));
 sky130_fd_sc_hd__and3_1 _4655_ (.A(\mem[29][27] ),
    .B(_1202_),
    .C(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__and3_1 _4656_ (.A(\mem[30][27] ),
    .B(_1232_),
    .C(_1013_),
    .X(_1323_));
 sky130_fd_sc_hd__a2111o_1 _4657_ (.A1(\mem[25][27] ),
    .A2(_0997_),
    .B1(_1320_),
    .C1(_1322_),
    .D1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__and3_1 _4658_ (.A(\mem[15][27] ),
    .B(_1107_),
    .C(_1235_),
    .X(_1325_));
 sky130_fd_sc_hd__buf_4 _4659_ (.A(_1021_),
    .X(_1326_));
 sky130_fd_sc_hd__and3_1 _4660_ (.A(\mem[24][27] ),
    .B(_1326_),
    .C(_1295_),
    .X(_1327_));
 sky130_fd_sc_hd__and3_1 _4661_ (.A(\mem[13][27] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1328_));
 sky130_fd_sc_hd__a2111o_1 _4662_ (.A1(\mem[10][27] ),
    .A2(_1017_),
    .B1(_1325_),
    .C1(_1327_),
    .D1(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__inv_2 _4663_ (.A(\mem[3][27] ),
    .Y(_1330_));
 sky130_fd_sc_hd__inv_2 _4664_ (.A(\mem[19][27] ),
    .Y(_1331_));
 sky130_fd_sc_hd__or3_1 _4665_ (.A(_1331_),
    .B(_1115_),
    .C(_1152_),
    .X(_1332_));
 sky130_fd_sc_hd__or3b_1 _4666_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][27] ),
    .X(_1333_));
 sky130_fd_sc_hd__or3b_1 _4667_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][27] ),
    .X(_1334_));
 sky130_fd_sc_hd__o2111ai_1 _4668_ (.A1(_1330_),
    .A2(_1035_),
    .B1(_1332_),
    .C1(_1333_),
    .D1(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__buf_4 _4669_ (.A(_1003_),
    .X(_1336_));
 sky130_fd_sc_hd__and3_1 _4670_ (.A(\mem[4][27] ),
    .B(_1336_),
    .C(_1275_),
    .X(_1337_));
 sky130_fd_sc_hd__buf_4 _4671_ (.A(_0995_),
    .X(_1338_));
 sky130_fd_sc_hd__buf_4 _4672_ (.A(_1058_),
    .X(_1339_));
 sky130_fd_sc_hd__and3_1 _4673_ (.A(\mem[22][27] ),
    .B(_1338_),
    .C(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__and3_1 _4674_ (.A(\mem[20][27] ),
    .B(_1061_),
    .C(_1063_),
    .X(_1341_));
 sky130_fd_sc_hd__a2111o_1 _4675_ (.A1(\mem[18][27] ),
    .A2(_1051_),
    .B1(_1337_),
    .C1(_1340_),
    .D1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__or4_1 _4676_ (.A(_1324_),
    .B(_1329_),
    .C(_1335_),
    .D(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__a22o_1 _4677_ (.A1(\mem[9][27] ),
    .A2(_1077_),
    .B1(_1079_),
    .B2(\mem[11][27] ),
    .X(_1344_));
 sky130_fd_sc_hd__a22o_1 _4678_ (.A1(\mem[27][27] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][27] ),
    .X(_1345_));
 sky130_fd_sc_hd__a32o_1 _4679_ (.A1(\mem[31][27] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][27] ),
    .X(_1346_));
 sky130_fd_sc_hd__a2111o_1 _4680_ (.A1(\mem[26][27] ),
    .A2(_1069_),
    .B1(_1344_),
    .C1(_1345_),
    .D1(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a22o_1 _4681_ (.A1(\mem[16][27] ),
    .A2(_1087_),
    .B1(_1089_),
    .B2(\mem[7][27] ),
    .X(_1348_));
 sky130_fd_sc_hd__a221o_1 _4682_ (.A1(\mem[8][27] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][27] ),
    .C1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a22o_1 _4683_ (.A1(\mem[21][27] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][27] ),
    .X(_1350_));
 sky130_fd_sc_hd__a221o_1 _4684_ (.A1(\mem[2][27] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][27] ),
    .C1(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__or4_4 _4685_ (.A(_1343_),
    .B(_1347_),
    .C(_1349_),
    .D(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _4686_ (.A(_1352_),
    .X(net101));
 sky130_fd_sc_hd__buf_6 _4687_ (.A(_0996_),
    .X(_1353_));
 sky130_fd_sc_hd__and3_1 _4688_ (.A(\mem[12][28] ),
    .B(_1319_),
    .C(_1260_),
    .X(_1354_));
 sky130_fd_sc_hd__and3_1 _4689_ (.A(\mem[29][28] ),
    .B(_1202_),
    .C(_1321_),
    .X(_1355_));
 sky130_fd_sc_hd__buf_4 _4690_ (.A(_1012_),
    .X(_1356_));
 sky130_fd_sc_hd__and3_1 _4691_ (.A(\mem[30][28] ),
    .B(_1232_),
    .C(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__a2111o_1 _4692_ (.A1(\mem[25][28] ),
    .A2(_1353_),
    .B1(_1354_),
    .C1(_1355_),
    .D1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__buf_4 _4693_ (.A(_1016_),
    .X(_1359_));
 sky130_fd_sc_hd__and3_1 _4694_ (.A(\mem[15][28] ),
    .B(_1107_),
    .C(_1235_),
    .X(_1360_));
 sky130_fd_sc_hd__and3_1 _4695_ (.A(\mem[24][28] ),
    .B(_1326_),
    .C(_1295_),
    .X(_1361_));
 sky130_fd_sc_hd__and3_1 _4696_ (.A(\mem[13][28] ),
    .B(_1147_),
    .C(_1110_),
    .X(_1362_));
 sky130_fd_sc_hd__a2111o_1 _4697_ (.A1(\mem[10][28] ),
    .A2(_1359_),
    .B1(_1360_),
    .C1(_1361_),
    .D1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__inv_2 _4698_ (.A(\mem[3][28] ),
    .Y(_1364_));
 sky130_fd_sc_hd__inv_2 _4699_ (.A(\mem[19][28] ),
    .Y(_1365_));
 sky130_fd_sc_hd__or3_1 _4700_ (.A(_1365_),
    .B(_1115_),
    .C(_1152_),
    .X(_1366_));
 sky130_fd_sc_hd__or3b_1 _4701_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][28] ),
    .X(_1367_));
 sky130_fd_sc_hd__or3b_1 _4702_ (.A(_1118_),
    .B(_1119_),
    .C_N(\mem[1][28] ),
    .X(_1368_));
 sky130_fd_sc_hd__o2111ai_1 _4703_ (.A1(_1364_),
    .A2(_1035_),
    .B1(_1366_),
    .C1(_1367_),
    .D1(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__buf_4 _4704_ (.A(_1050_),
    .X(_1370_));
 sky130_fd_sc_hd__and3_1 _4705_ (.A(\mem[4][28] ),
    .B(_1336_),
    .C(_1275_),
    .X(_1371_));
 sky130_fd_sc_hd__and3_1 _4706_ (.A(\mem[22][28] ),
    .B(_1338_),
    .C(_1339_),
    .X(_1372_));
 sky130_fd_sc_hd__buf_4 _4707_ (.A(_1054_),
    .X(_1373_));
 sky130_fd_sc_hd__buf_4 _4708_ (.A(_1062_),
    .X(_1374_));
 sky130_fd_sc_hd__and3_1 _4709_ (.A(\mem[20][28] ),
    .B(_1373_),
    .C(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__a2111o_1 _4710_ (.A1(\mem[18][28] ),
    .A2(_1370_),
    .B1(_1371_),
    .C1(_1372_),
    .D1(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__or4_1 _4711_ (.A(_1358_),
    .B(_1363_),
    .C(_1369_),
    .D(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__buf_6 _4712_ (.A(_1076_),
    .X(_1378_));
 sky130_fd_sc_hd__a22o_1 _4713_ (.A1(\mem[9][28] ),
    .A2(_1378_),
    .B1(_1079_),
    .B2(\mem[11][28] ),
    .X(_1379_));
 sky130_fd_sc_hd__a22o_1 _4714_ (.A1(\mem[27][28] ),
    .A2(_1128_),
    .B1(_1129_),
    .B2(\mem[28][28] ),
    .X(_1380_));
 sky130_fd_sc_hd__a32o_1 _4715_ (.A1(\mem[31][28] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(\mem[14][28] ),
    .X(_1381_));
 sky130_fd_sc_hd__a2111o_1 _4716_ (.A1(\mem[26][28] ),
    .A2(_1069_),
    .B1(_1379_),
    .C1(_1380_),
    .D1(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__buf_6 _4717_ (.A(_1086_),
    .X(_1383_));
 sky130_fd_sc_hd__buf_6 _4718_ (.A(_1088_),
    .X(_1384_));
 sky130_fd_sc_hd__a22o_1 _4719_ (.A1(\mem[16][28] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][28] ),
    .X(_1385_));
 sky130_fd_sc_hd__a221o_1 _4720_ (.A1(\mem[8][28] ),
    .A2(_1083_),
    .B1(_1085_),
    .B2(\mem[6][28] ),
    .C1(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__a22o_1 _4721_ (.A1(\mem[21][28] ),
    .A2(_1097_),
    .B1(_1099_),
    .B2(\mem[17][28] ),
    .X(_1387_));
 sky130_fd_sc_hd__a221o_1 _4722_ (.A1(\mem[2][28] ),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\mem[23][28] ),
    .C1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__or4_4 _4723_ (.A(_1377_),
    .B(_1382_),
    .C(_1386_),
    .D(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__buf_2 _4724_ (.A(_1389_),
    .X(net102));
 sky130_fd_sc_hd__and3_1 _4725_ (.A(\mem[12][29] ),
    .B(_1319_),
    .C(_1260_),
    .X(_1390_));
 sky130_fd_sc_hd__and3_1 _4726_ (.A(\mem[29][29] ),
    .B(_1202_),
    .C(_1321_),
    .X(_1391_));
 sky130_fd_sc_hd__and3_1 _4727_ (.A(\mem[30][29] ),
    .B(_1232_),
    .C(_1356_),
    .X(_1392_));
 sky130_fd_sc_hd__a2111o_1 _4728_ (.A1(\mem[25][29] ),
    .A2(_1353_),
    .B1(_1390_),
    .C1(_1391_),
    .D1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__and3_1 _4729_ (.A(\mem[15][29] ),
    .B(_1107_),
    .C(_1235_),
    .X(_1394_));
 sky130_fd_sc_hd__and3_1 _4730_ (.A(\mem[24][29] ),
    .B(_1326_),
    .C(_1295_),
    .X(_1395_));
 sky130_fd_sc_hd__buf_4 _4731_ (.A(_1007_),
    .X(_1396_));
 sky130_fd_sc_hd__and3_1 _4732_ (.A(\mem[13][29] ),
    .B(_1147_),
    .C(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__a2111o_1 _4733_ (.A1(\mem[10][29] ),
    .A2(_1359_),
    .B1(_1394_),
    .C1(_1395_),
    .D1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__inv_2 _4734_ (.A(\mem[3][29] ),
    .Y(_1399_));
 sky130_fd_sc_hd__buf_4 _4735_ (.A(_1034_),
    .X(_1400_));
 sky130_fd_sc_hd__inv_2 _4736_ (.A(\mem[19][29] ),
    .Y(_1401_));
 sky130_fd_sc_hd__or3_1 _4737_ (.A(_1401_),
    .B(_1115_),
    .C(_1152_),
    .X(_1402_));
 sky130_fd_sc_hd__or3b_1 _4738_ (.A(_1039_),
    .B(_1041_),
    .C_N(\mem[5][29] ),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_4 _4739_ (.A(_1037_),
    .X(_1404_));
 sky130_fd_sc_hd__or3b_1 _4740_ (.A(_1118_),
    .B(_1404_),
    .C_N(\mem[1][29] ),
    .X(_1405_));
 sky130_fd_sc_hd__o2111ai_1 _4741_ (.A1(_1399_),
    .A2(_1400_),
    .B1(_1402_),
    .C1(_1403_),
    .D1(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__and3_1 _4742_ (.A(\mem[4][29] ),
    .B(_1336_),
    .C(_1275_),
    .X(_1407_));
 sky130_fd_sc_hd__and3_1 _4743_ (.A(\mem[22][29] ),
    .B(_1338_),
    .C(_1339_),
    .X(_1408_));
 sky130_fd_sc_hd__and3_1 _4744_ (.A(\mem[20][29] ),
    .B(_1373_),
    .C(_1374_),
    .X(_1409_));
 sky130_fd_sc_hd__a2111o_1 _4745_ (.A1(\mem[18][29] ),
    .A2(_1370_),
    .B1(_1407_),
    .C1(_1408_),
    .D1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__or4_1 _4746_ (.A(_1393_),
    .B(_1398_),
    .C(_1406_),
    .D(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__buf_6 _4747_ (.A(_1068_),
    .X(_1412_));
 sky130_fd_sc_hd__buf_6 _4748_ (.A(_1078_),
    .X(_1413_));
 sky130_fd_sc_hd__a22o_1 _4749_ (.A1(\mem[9][29] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][29] ),
    .X(_1414_));
 sky130_fd_sc_hd__buf_6 _4750_ (.A(_1070_),
    .X(_1415_));
 sky130_fd_sc_hd__a22o_1 _4751_ (.A1(\mem[27][29] ),
    .A2(_1415_),
    .B1(_1129_),
    .B2(\mem[28][29] ),
    .X(_1416_));
 sky130_fd_sc_hd__buf_6 _4752_ (.A(_1074_),
    .X(_1417_));
 sky130_fd_sc_hd__a32o_1 _4753_ (.A1(\mem[31][29] ),
    .A2(_1193_),
    .A3(_1132_),
    .B1(_1417_),
    .B2(\mem[14][29] ),
    .X(_1418_));
 sky130_fd_sc_hd__a2111o_1 _4754_ (.A1(\mem[26][29] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1416_),
    .D1(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_8 _4755_ (.A(_1082_),
    .X(_1420_));
 sky130_fd_sc_hd__buf_6 _4756_ (.A(_1084_),
    .X(_1421_));
 sky130_fd_sc_hd__a22o_1 _4757_ (.A1(\mem[16][29] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][29] ),
    .X(_1422_));
 sky130_fd_sc_hd__a221o_1 _4758_ (.A1(\mem[8][29] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][29] ),
    .C1(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_8 _4759_ (.A(_1092_),
    .X(_1424_));
 sky130_fd_sc_hd__buf_4 _4760_ (.A(_1094_),
    .X(_1425_));
 sky130_fd_sc_hd__buf_6 _4761_ (.A(_1096_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_8 _4762_ (.A(_1098_),
    .X(_1427_));
 sky130_fd_sc_hd__a22o_1 _4763_ (.A1(\mem[21][29] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][29] ),
    .X(_1428_));
 sky130_fd_sc_hd__a221o_1 _4764_ (.A1(\mem[2][29] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][29] ),
    .C1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__or4_4 _4765_ (.A(_1411_),
    .B(_1419_),
    .C(_1423_),
    .D(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_4 _4766_ (.A(_1430_),
    .X(net103));
 sky130_fd_sc_hd__and3_1 _4767_ (.A(\mem[12][30] ),
    .B(_1319_),
    .C(_1260_),
    .X(_1431_));
 sky130_fd_sc_hd__and3_1 _4768_ (.A(\mem[29][30] ),
    .B(_1202_),
    .C(_1321_),
    .X(_1432_));
 sky130_fd_sc_hd__and3_1 _4769_ (.A(\mem[30][30] ),
    .B(_1232_),
    .C(_1356_),
    .X(_1433_));
 sky130_fd_sc_hd__a2111o_1 _4770_ (.A1(\mem[25][30] ),
    .A2(_1353_),
    .B1(_1431_),
    .C1(_1432_),
    .D1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_4 _4771_ (.A(_1018_),
    .X(_1435_));
 sky130_fd_sc_hd__and3_1 _4772_ (.A(\mem[15][30] ),
    .B(_1435_),
    .C(_1235_),
    .X(_1436_));
 sky130_fd_sc_hd__and3_1 _4773_ (.A(\mem[24][30] ),
    .B(_1326_),
    .C(_1295_),
    .X(_1437_));
 sky130_fd_sc_hd__and3_1 _4774_ (.A(\mem[13][30] ),
    .B(_1147_),
    .C(_1396_),
    .X(_1438_));
 sky130_fd_sc_hd__a2111o_1 _4775_ (.A1(\mem[10][30] ),
    .A2(_1359_),
    .B1(_1436_),
    .C1(_1437_),
    .D1(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__inv_2 _4776_ (.A(\mem[3][30] ),
    .Y(_1440_));
 sky130_fd_sc_hd__inv_2 _4777_ (.A(\mem[19][30] ),
    .Y(_1441_));
 sky130_fd_sc_hd__or3_1 _4778_ (.A(_1441_),
    .B(_1115_),
    .C(_1152_),
    .X(_1442_));
 sky130_fd_sc_hd__buf_2 _4779_ (.A(_1040_),
    .X(_1443_));
 sky130_fd_sc_hd__or3b_1 _4780_ (.A(_1039_),
    .B(_1443_),
    .C_N(\mem[5][30] ),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_4 _4781_ (.A(_1010_),
    .X(_1445_));
 sky130_fd_sc_hd__or3b_1 _4782_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][30] ),
    .X(_1446_));
 sky130_fd_sc_hd__o2111ai_1 _4783_ (.A1(_1440_),
    .A2(_1400_),
    .B1(_1442_),
    .C1(_1444_),
    .D1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__and3_1 _4784_ (.A(\mem[4][30] ),
    .B(_1336_),
    .C(_1275_),
    .X(_1448_));
 sky130_fd_sc_hd__and3_1 _4785_ (.A(\mem[22][30] ),
    .B(_1338_),
    .C(_1339_),
    .X(_1449_));
 sky130_fd_sc_hd__and3_1 _4786_ (.A(\mem[20][30] ),
    .B(_1373_),
    .C(_1374_),
    .X(_1450_));
 sky130_fd_sc_hd__a2111o_1 _4787_ (.A1(\mem[18][30] ),
    .A2(_1370_),
    .B1(_1448_),
    .C1(_1449_),
    .D1(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__or4_1 _4788_ (.A(_1434_),
    .B(_1439_),
    .C(_1447_),
    .D(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__a22o_1 _4789_ (.A1(\mem[9][30] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][30] ),
    .X(_1453_));
 sky130_fd_sc_hd__buf_6 _4790_ (.A(_1071_),
    .X(_1454_));
 sky130_fd_sc_hd__a22o_1 _4791_ (.A1(\mem[27][30] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][30] ),
    .X(_1455_));
 sky130_fd_sc_hd__buf_6 _4792_ (.A(_1028_),
    .X(_1456_));
 sky130_fd_sc_hd__a32o_1 _4793_ (.A1(\mem[31][30] ),
    .A2(_1193_),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][30] ),
    .X(_1457_));
 sky130_fd_sc_hd__a2111o_1 _4794_ (.A1(\mem[26][30] ),
    .A2(_1412_),
    .B1(_1453_),
    .C1(_1455_),
    .D1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__a22o_1 _4795_ (.A1(\mem[16][30] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][30] ),
    .X(_1459_));
 sky130_fd_sc_hd__a221o_1 _4796_ (.A1(\mem[8][30] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][30] ),
    .C1(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a22o_1 _4797_ (.A1(\mem[21][30] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][30] ),
    .X(_1461_));
 sky130_fd_sc_hd__a221o_1 _4798_ (.A1(\mem[2][30] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][30] ),
    .C1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__or4_4 _4799_ (.A(_1452_),
    .B(_1458_),
    .C(_1460_),
    .D(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _4800_ (.A(_1463_),
    .X(net105));
 sky130_fd_sc_hd__and3_1 _4801_ (.A(\mem[12][31] ),
    .B(_1319_),
    .C(_1260_),
    .X(_1464_));
 sky130_fd_sc_hd__and3_1 _4802_ (.A(\mem[29][31] ),
    .B(_1202_),
    .C(_1321_),
    .X(_1465_));
 sky130_fd_sc_hd__and3_1 _4803_ (.A(\mem[30][31] ),
    .B(_1232_),
    .C(_1356_),
    .X(_1466_));
 sky130_fd_sc_hd__a2111o_1 _4804_ (.A1(\mem[25][31] ),
    .A2(_1353_),
    .B1(_1464_),
    .C1(_1465_),
    .D1(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__and3_1 _4805_ (.A(\mem[15][31] ),
    .B(_1435_),
    .C(_1235_),
    .X(_1468_));
 sky130_fd_sc_hd__and3_1 _4806_ (.A(\mem[24][31] ),
    .B(_1326_),
    .C(_1295_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_4 _4807_ (.A(_1044_),
    .X(_1470_));
 sky130_fd_sc_hd__and3_1 _4808_ (.A(\mem[13][31] ),
    .B(_1470_),
    .C(_1396_),
    .X(_1471_));
 sky130_fd_sc_hd__a2111o_1 _4809_ (.A1(\mem[10][31] ),
    .A2(_1359_),
    .B1(_1468_),
    .C1(_1469_),
    .D1(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__inv_2 _4810_ (.A(\mem[3][31] ),
    .Y(_1473_));
 sky130_fd_sc_hd__inv_2 _4811_ (.A(\mem[19][31] ),
    .Y(_1474_));
 sky130_fd_sc_hd__or3_1 _4812_ (.A(_1474_),
    .B(_1115_),
    .C(_1152_),
    .X(_1475_));
 sky130_fd_sc_hd__or3b_1 _4813_ (.A(_1039_),
    .B(_1443_),
    .C_N(\mem[5][31] ),
    .X(_1476_));
 sky130_fd_sc_hd__or3b_1 _4814_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][31] ),
    .X(_1477_));
 sky130_fd_sc_hd__o2111ai_1 _4815_ (.A1(_1473_),
    .A2(_1400_),
    .B1(_1475_),
    .C1(_1476_),
    .D1(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__and3_1 _4816_ (.A(\mem[4][31] ),
    .B(_1336_),
    .C(_1275_),
    .X(_1479_));
 sky130_fd_sc_hd__and3_1 _4817_ (.A(\mem[22][31] ),
    .B(_1338_),
    .C(_1339_),
    .X(_1480_));
 sky130_fd_sc_hd__and3_1 _4818_ (.A(\mem[20][31] ),
    .B(_1373_),
    .C(_1374_),
    .X(_1481_));
 sky130_fd_sc_hd__a2111o_1 _4819_ (.A1(\mem[18][31] ),
    .A2(_1370_),
    .B1(_1479_),
    .C1(_1480_),
    .D1(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__or4_1 _4820_ (.A(_1467_),
    .B(_1472_),
    .C(_1478_),
    .D(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__a22o_1 _4821_ (.A1(\mem[9][31] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][31] ),
    .X(_1484_));
 sky130_fd_sc_hd__a22o_1 _4822_ (.A1(\mem[27][31] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][31] ),
    .X(_1485_));
 sky130_fd_sc_hd__a32o_1 _4823_ (.A1(\mem[31][31] ),
    .A2(_1193_),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][31] ),
    .X(_1486_));
 sky130_fd_sc_hd__a2111o_1 _4824_ (.A1(\mem[26][31] ),
    .A2(_1412_),
    .B1(_1484_),
    .C1(_1485_),
    .D1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__a22o_1 _4825_ (.A1(\mem[16][31] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][31] ),
    .X(_1488_));
 sky130_fd_sc_hd__a221o_1 _4826_ (.A1(\mem[8][31] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][31] ),
    .C1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__a22o_1 _4827_ (.A1(\mem[21][31] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][31] ),
    .X(_1490_));
 sky130_fd_sc_hd__a221o_1 _4828_ (.A1(\mem[2][31] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][31] ),
    .C1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__or4_4 _4829_ (.A(_1483_),
    .B(_1487_),
    .C(_1489_),
    .D(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_4 _4830_ (.A(_1492_),
    .X(net106));
 sky130_fd_sc_hd__inv_2 _4831_ (.A(net5),
    .Y(_1493_));
 sky130_fd_sc_hd__clkbuf_4 _4832_ (.A(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_4 _4833_ (.A(net1),
    .X(_1495_));
 sky130_fd_sc_hd__buf_2 _4834_ (.A(net2),
    .X(_1496_));
 sky130_fd_sc_hd__and4b_2 _4835_ (.A_N(net3),
    .B(net4),
    .C(_1495_),
    .D(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__and2_2 _4836_ (.A(_1494_),
    .B(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__buf_2 _4837_ (.A(net5),
    .X(_1499_));
 sky130_fd_sc_hd__and4_2 _4838_ (.A(net2),
    .B(net1),
    .C(net4),
    .D(net3),
    .X(_1500_));
 sky130_fd_sc_hd__and2_2 _4839_ (.A(_1499_),
    .B(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__a22o_1 _4840_ (.A1(\mem[11][0] ),
    .A2(_1498_),
    .B1(_1501_),
    .B2(\mem[31][0] ),
    .X(_1502_));
 sky130_fd_sc_hd__nor2_1 _4841_ (.A(net4),
    .B(net3),
    .Y(_1503_));
 sky130_fd_sc_hd__clkbuf_4 _4842_ (.A(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_4 _4843_ (.A(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__and3b_2 _4844_ (.A_N(net1),
    .B(net2),
    .C(net5),
    .X(_1506_));
 sky130_fd_sc_hd__buf_2 _4845_ (.A(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_4 _4846_ (.A(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__and2_2 _4847_ (.A(net4),
    .B(net3),
    .X(_1509_));
 sky130_fd_sc_hd__nor2_1 _4848_ (.A(_1496_),
    .B(_1495_),
    .Y(_1510_));
 sky130_fd_sc_hd__and3_2 _4849_ (.A(_1493_),
    .B(_1509_),
    .C(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__buf_4 _4850_ (.A(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__a32o_1 _4851_ (.A1(\mem[18][0] ),
    .A2(_1505_),
    .A3(_1508_),
    .B1(\mem[12][0] ),
    .B2(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__buf_4 _4852_ (.A(_1499_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_4 _4853_ (.A(_1497_),
    .X(_1515_));
 sky130_fd_sc_hd__buf_2 _4854_ (.A(net3),
    .X(_1516_));
 sky130_fd_sc_hd__buf_2 _4855_ (.A(net4),
    .X(_1517_));
 sky130_fd_sc_hd__and2b_1 _4856_ (.A_N(_1516_),
    .B(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__buf_2 _4857_ (.A(net5),
    .X(_1519_));
 sky130_fd_sc_hd__and4b_2 _4858_ (.A_N(_1496_),
    .B(_1495_),
    .C(_1518_),
    .D(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__a32o_1 _4859_ (.A1(_1514_),
    .A2(\mem[27][0] ),
    .A3(_1515_),
    .B1(_1520_),
    .B2(\mem[25][0] ),
    .X(_1521_));
 sky130_fd_sc_hd__nor4b_4 _4860_ (.A(_1496_),
    .B(_1495_),
    .C(net3),
    .D_N(net4),
    .Y(_1522_));
 sky130_fd_sc_hd__clkbuf_4 _4861_ (.A(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__nor3b_4 _4862_ (.A(net5),
    .B(_1495_),
    .C_N(_1496_),
    .Y(_1524_));
 sky130_fd_sc_hd__and2_2 _4863_ (.A(_1509_),
    .B(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__a32o_1 _4864_ (.A1(_1514_),
    .A2(\mem[24][0] ),
    .A3(_1523_),
    .B1(_1525_),
    .B2(\mem[14][0] ),
    .X(_1526_));
 sky130_fd_sc_hd__or4_1 _4865_ (.A(_1502_),
    .B(_1513_),
    .C(_1521_),
    .D(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__or3b_2 _4866_ (.A(_1517_),
    .B(_1516_),
    .C_N(net5),
    .X(_1528_));
 sky130_fd_sc_hd__or2b_1 _4867_ (.A(_1496_),
    .B_N(_1495_),
    .X(_1529_));
 sky130_fd_sc_hd__nor2_2 _4868_ (.A(_1528_),
    .B(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__buf_4 _4869_ (.A(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_4 _4870_ (.A(_1493_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_4 _4871_ (.A(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_4 _4872_ (.A(_1500_),
    .X(_1534_));
 sky130_fd_sc_hd__and3_1 _4873_ (.A(_1533_),
    .B(\mem[15][0] ),
    .C(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__buf_4 _4874_ (.A(_1517_),
    .X(_1536_));
 sky130_fd_sc_hd__buf_4 _4875_ (.A(_1516_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_4 _4876_ (.A(_1524_),
    .X(_1538_));
 sky130_fd_sc_hd__and3b_2 _4877_ (.A_N(_1536_),
    .B(_1537_),
    .C(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__or4b_2 _4878_ (.A(net2),
    .B(net1),
    .C(net4),
    .D_N(net3),
    .X(_1540_));
 sky130_fd_sc_hd__nor2_4 _4879_ (.A(_1532_),
    .B(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__buf_4 _4880_ (.A(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_4 _4881_ (.A(_1509_),
    .X(_1543_));
 sky130_fd_sc_hd__and4_1 _4882_ (.A(_1514_),
    .B(\mem[28][0] ),
    .C(_1543_),
    .D(_1510_),
    .X(_1544_));
 sky130_fd_sc_hd__a221o_1 _4883_ (.A1(\mem[6][0] ),
    .A2(_1539_),
    .B1(_1542_),
    .B2(\mem[20][0] ),
    .C1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__and3_2 _4884_ (.A(_1499_),
    .B(_1510_),
    .C(_1504_),
    .X(_1546_));
 sky130_fd_sc_hd__buf_4 _4885_ (.A(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__or3_1 _4886_ (.A(net5),
    .B(net4),
    .C(net3),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_2 _4887_ (.A(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__nor2_2 _4888_ (.A(_1529_),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__clkbuf_4 _4889_ (.A(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__a22o_1 _4890_ (.A1(\mem[16][0] ),
    .A2(_1547_),
    .B1(_1551_),
    .B2(\mem[1][0] ),
    .X(_1552_));
 sky130_fd_sc_hd__a2111o_1 _4891_ (.A1(\mem[17][0] ),
    .A2(_1531_),
    .B1(_1535_),
    .C1(_1545_),
    .D1(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__nor2_4 _4892_ (.A(_1514_),
    .B(_1540_),
    .Y(_1554_));
 sky130_fd_sc_hd__inv_2 _4893_ (.A(\mem[21][0] ),
    .Y(_1555_));
 sky130_fd_sc_hd__or4bb_4 _4894_ (.A(_1496_),
    .B(net4),
    .C_N(net3),
    .D_N(_1495_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_4 _4895_ (.A(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__nor3_1 _4896_ (.A(_1533_),
    .B(_1555_),
    .C(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__and3_1 _4897_ (.A(\mem[2][0] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1559_));
 sky130_fd_sc_hd__nand4b_4 _4898_ (.A_N(_1496_),
    .B(_1495_),
    .C(_1517_),
    .D(_1516_),
    .Y(_1560_));
 sky130_fd_sc_hd__clkbuf_4 _4899_ (.A(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__and3b_1 _4900_ (.A_N(_1561_),
    .B(_1533_),
    .C(\mem[13][0] ),
    .X(_1562_));
 sky130_fd_sc_hd__a2111oi_1 _4901_ (.A1(\mem[4][0] ),
    .A2(_1554_),
    .B1(_1558_),
    .C1(_1559_),
    .D1(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__and4b_2 _4902_ (.A_N(_1517_),
    .B(_1516_),
    .C(_1496_),
    .D(_1495_),
    .X(_1564_));
 sky130_fd_sc_hd__and2_2 _4903_ (.A(_1494_),
    .B(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__buf_4 _4904_ (.A(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__and3_1 _4905_ (.A(\mem[30][0] ),
    .B(_1543_),
    .C(_1508_),
    .X(_1567_));
 sky130_fd_sc_hd__and3b_1 _4906_ (.A_N(_1557_),
    .B(_1533_),
    .C(\mem[5][0] ),
    .X(_1568_));
 sky130_fd_sc_hd__and3_1 _4907_ (.A(\mem[10][0] ),
    .B(_1518_),
    .C(_1538_),
    .X(_1569_));
 sky130_fd_sc_hd__a2111oi_1 _4908_ (.A1(\mem[7][0] ),
    .A2(_1566_),
    .B1(_1567_),
    .C1(_1568_),
    .D1(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__and3b_2 _4909_ (.A_N(_1529_),
    .B(_1494_),
    .C(_1518_),
    .X(_1571_));
 sky130_fd_sc_hd__buf_4 _4910_ (.A(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_4 _4911_ (.A(_1564_),
    .X(_1573_));
 sky130_fd_sc_hd__and3_1 _4912_ (.A(_1514_),
    .B(\mem[23][0] ),
    .C(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__inv_2 _4913_ (.A(\mem[29][0] ),
    .Y(_1575_));
 sky130_fd_sc_hd__nor3_1 _4914_ (.A(_1533_),
    .B(_1575_),
    .C(_1561_),
    .Y(_1576_));
 sky130_fd_sc_hd__and3_1 _4915_ (.A(\mem[26][0] ),
    .B(_1518_),
    .C(_1508_),
    .X(_1577_));
 sky130_fd_sc_hd__a2111oi_1 _4916_ (.A1(\mem[9][0] ),
    .A2(_1572_),
    .B1(_1574_),
    .C1(_1576_),
    .D1(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_2 _4917_ (.A(_1496_),
    .B(_1495_),
    .Y(_1579_));
 sky130_fd_sc_hd__nor2_4 _4918_ (.A(_1579_),
    .B(_1528_),
    .Y(_1580_));
 sky130_fd_sc_hd__buf_4 _4919_ (.A(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__and4b_1 _4920_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][0] ),
    .D(_1508_),
    .X(_1582_));
 sky130_fd_sc_hd__and3_1 _4921_ (.A(_1533_),
    .B(\mem[8][0] ),
    .C(_1523_),
    .X(_1583_));
 sky130_fd_sc_hd__buf_4 _4922_ (.A(_1579_),
    .X(_1584_));
 sky130_fd_sc_hd__and4b_1 _4923_ (.A_N(_1584_),
    .B(_1533_),
    .C(\mem[3][0] ),
    .D(_1505_),
    .X(_1585_));
 sky130_fd_sc_hd__a2111oi_1 _4924_ (.A1(\mem[19][0] ),
    .A2(_1581_),
    .B1(_1582_),
    .C1(_1583_),
    .D1(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__and4_1 _4925_ (.A(_1563_),
    .B(_1570_),
    .C(_1578_),
    .D(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__or3b_4 _4926_ (.A(_1527_),
    .B(_1553_),
    .C_N(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _4927_ (.A(_1588_),
    .X(net50));
 sky130_fd_sc_hd__buf_4 _4928_ (.A(_1519_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_4 _4929_ (.A(_1522_),
    .X(_1590_));
 sky130_fd_sc_hd__and3_1 _4930_ (.A(_1589_),
    .B(\mem[24][1] ),
    .C(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__buf_4 _4931_ (.A(_1506_),
    .X(_1592_));
 sky130_fd_sc_hd__and3_1 _4932_ (.A(\mem[30][1] ),
    .B(_1543_),
    .C(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_4 _4933_ (.A(_1519_),
    .X(_1594_));
 sky130_fd_sc_hd__and3_1 _4934_ (.A(_1594_),
    .B(\mem[27][1] ),
    .C(_1515_),
    .X(_1595_));
 sky130_fd_sc_hd__a2111o_1 _4935_ (.A1(\mem[12][1] ),
    .A2(_1512_),
    .B1(_1591_),
    .C1(_1593_),
    .D1(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__and2_1 _4936_ (.A(_1518_),
    .B(_1524_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_4 _4937_ (.A(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__buf_4 _4938_ (.A(_1532_),
    .X(_1599_));
 sky130_fd_sc_hd__and3_1 _4939_ (.A(_1599_),
    .B(\mem[15][1] ),
    .C(_1534_),
    .X(_1600_));
 sky130_fd_sc_hd__buf_4 _4940_ (.A(_1560_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_4 _4941_ (.A(_1532_),
    .X(_1602_));
 sky130_fd_sc_hd__and3b_1 _4942_ (.A_N(_1601_),
    .B(_1602_),
    .C(\mem[13][1] ),
    .X(_1603_));
 sky130_fd_sc_hd__and3_1 _4943_ (.A(_1533_),
    .B(\mem[8][1] ),
    .C(_1523_),
    .X(_1604_));
 sky130_fd_sc_hd__a2111o_1 _4944_ (.A1(\mem[10][1] ),
    .A2(_1598_),
    .B1(_1600_),
    .C1(_1603_),
    .D1(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__inv_2 _4945_ (.A(\mem[3][1] ),
    .Y(_1606_));
 sky130_fd_sc_hd__buf_4 _4946_ (.A(_1579_),
    .X(_1607_));
 sky130_fd_sc_hd__buf_4 _4947_ (.A(_1549_),
    .X(_1608_));
 sky130_fd_sc_hd__nor3_1 _4948_ (.A(_1606_),
    .B(_1607_),
    .C(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__buf_4 _4949_ (.A(_1506_),
    .X(_1610_));
 sky130_fd_sc_hd__and4b_1 _4950_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][1] ),
    .D(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__buf_4 _4951_ (.A(_1556_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_4 _4952_ (.A(_1532_),
    .X(_1613_));
 sky130_fd_sc_hd__and3b_1 _4953_ (.A_N(_1612_),
    .B(_1613_),
    .C(\mem[5][1] ),
    .X(_1614_));
 sky130_fd_sc_hd__a2111o_1 _4954_ (.A1(\mem[1][1] ),
    .A2(_1551_),
    .B1(_1609_),
    .C1(_1611_),
    .D1(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__buf_4 _4955_ (.A(_1504_),
    .X(_1616_));
 sky130_fd_sc_hd__and3_1 _4956_ (.A(\mem[18][1] ),
    .B(_1616_),
    .C(_1508_),
    .X(_1617_));
 sky130_fd_sc_hd__and3_1 _4957_ (.A(\mem[2][1] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1618_));
 sky130_fd_sc_hd__buf_4 _4958_ (.A(_1519_),
    .X(_1619_));
 sky130_fd_sc_hd__and3_1 _4959_ (.A(_1619_),
    .B(\mem[23][1] ),
    .C(_1573_),
    .X(_1620_));
 sky130_fd_sc_hd__a2111o_1 _4960_ (.A1(\mem[20][1] ),
    .A2(_1542_),
    .B1(_1617_),
    .C1(_1618_),
    .D1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__or4_1 _4961_ (.A(_1596_),
    .B(_1605_),
    .C(_1615_),
    .D(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__and2_2 _4962_ (.A(_1518_),
    .B(_1508_),
    .X(_1623_));
 sky130_fd_sc_hd__buf_4 _4963_ (.A(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__a22o_1 _4964_ (.A1(\mem[7][1] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][1] ),
    .X(_1625_));
 sky130_fd_sc_hd__buf_4 _4965_ (.A(_1501_),
    .X(_1626_));
 sky130_fd_sc_hd__buf_4 _4966_ (.A(_1520_),
    .X(_1627_));
 sky130_fd_sc_hd__a22o_1 _4967_ (.A1(\mem[31][1] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][1] ),
    .X(_1628_));
 sky130_fd_sc_hd__buf_4 _4968_ (.A(_1498_),
    .X(_1629_));
 sky130_fd_sc_hd__buf_4 _4969_ (.A(_1525_),
    .X(_1630_));
 sky130_fd_sc_hd__a22o_1 _4970_ (.A1(\mem[11][1] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][1] ),
    .X(_1631_));
 sky130_fd_sc_hd__a2111o_1 _4971_ (.A1(\mem[26][1] ),
    .A2(_1624_),
    .B1(_1625_),
    .C1(_1628_),
    .D1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__buf_4 _4972_ (.A(_1539_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_8 _4973_ (.A(_1554_),
    .X(_1634_));
 sky130_fd_sc_hd__a22o_1 _4974_ (.A1(\mem[16][1] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][1] ),
    .X(_1635_));
 sky130_fd_sc_hd__a221o_1 _4975_ (.A1(\mem[6][1] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][1] ),
    .C1(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__nor2_2 _4976_ (.A(_1533_),
    .B(_1557_),
    .Y(_1637_));
 sky130_fd_sc_hd__buf_4 _4977_ (.A(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__and3_2 _4978_ (.A(_1499_),
    .B(_1509_),
    .C(_1510_),
    .X(_1639_));
 sky130_fd_sc_hd__buf_4 _4979_ (.A(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__nor2_2 _4980_ (.A(_1533_),
    .B(_1601_),
    .Y(_1641_));
 sky130_fd_sc_hd__buf_4 _4981_ (.A(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__a22o_1 _4982_ (.A1(\mem[28][1] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][1] ),
    .X(_1643_));
 sky130_fd_sc_hd__a221o_1 _4983_ (.A1(\mem[17][1] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][1] ),
    .C1(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__or4_4 _4984_ (.A(_1622_),
    .B(_1632_),
    .C(_1636_),
    .D(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _4985_ (.A(_1645_),
    .X(net61));
 sky130_fd_sc_hd__and3_1 _4986_ (.A(_1589_),
    .B(\mem[24][2] ),
    .C(_1590_),
    .X(_1646_));
 sky130_fd_sc_hd__and3_1 _4987_ (.A(\mem[30][2] ),
    .B(_1543_),
    .C(_1592_),
    .X(_1647_));
 sky130_fd_sc_hd__and3_1 _4988_ (.A(_1594_),
    .B(\mem[27][2] ),
    .C(_1515_),
    .X(_1648_));
 sky130_fd_sc_hd__a2111o_1 _4989_ (.A1(\mem[12][2] ),
    .A2(_1512_),
    .B1(_1646_),
    .C1(_1647_),
    .D1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__and3_1 _4990_ (.A(_1599_),
    .B(\mem[15][2] ),
    .C(_1534_),
    .X(_1650_));
 sky130_fd_sc_hd__and3b_1 _4991_ (.A_N(_1601_),
    .B(_1602_),
    .C(\mem[13][2] ),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_4 _4992_ (.A(_1532_),
    .X(_1652_));
 sky130_fd_sc_hd__and3_1 _4993_ (.A(_1652_),
    .B(\mem[8][2] ),
    .C(_1523_),
    .X(_1653_));
 sky130_fd_sc_hd__a2111o_1 _4994_ (.A1(\mem[10][2] ),
    .A2(_1598_),
    .B1(_1650_),
    .C1(_1651_),
    .D1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_4 _4995_ (.A(_1517_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_4 _4996_ (.A(_1516_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_4 _4997_ (.A(_1506_),
    .X(_1657_));
 sky130_fd_sc_hd__and4b_1 _4998_ (.A_N(_1655_),
    .B(_1656_),
    .C(\mem[22][2] ),
    .D(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__inv_2 _4999_ (.A(\mem[3][2] ),
    .Y(_1659_));
 sky130_fd_sc_hd__buf_4 _5000_ (.A(_1549_),
    .X(_1660_));
 sky130_fd_sc_hd__nor3_1 _5001_ (.A(_1659_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__and3b_1 _5002_ (.A_N(_1612_),
    .B(_1613_),
    .C(\mem[5][2] ),
    .X(_1662_));
 sky130_fd_sc_hd__a2111o_1 _5003_ (.A1(\mem[1][2] ),
    .A2(_1551_),
    .B1(_1658_),
    .C1(_1661_),
    .D1(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__and3_1 _5004_ (.A(\mem[18][2] ),
    .B(_1616_),
    .C(_1508_),
    .X(_1664_));
 sky130_fd_sc_hd__and3_1 _5005_ (.A(\mem[2][2] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1665_));
 sky130_fd_sc_hd__and3_1 _5006_ (.A(_1619_),
    .B(\mem[23][2] ),
    .C(_1573_),
    .X(_1666_));
 sky130_fd_sc_hd__a2111o_1 _5007_ (.A1(\mem[20][2] ),
    .A2(_1542_),
    .B1(_1664_),
    .C1(_1665_),
    .D1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__or4_1 _5008_ (.A(_1649_),
    .B(_1654_),
    .C(_1663_),
    .D(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__a22o_1 _5009_ (.A1(\mem[7][2] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][2] ),
    .X(_1669_));
 sky130_fd_sc_hd__a22o_1 _5010_ (.A1(\mem[31][2] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][2] ),
    .X(_1670_));
 sky130_fd_sc_hd__a22o_1 _5011_ (.A1(\mem[11][2] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][2] ),
    .X(_1671_));
 sky130_fd_sc_hd__a2111o_1 _5012_ (.A1(\mem[26][2] ),
    .A2(_1624_),
    .B1(_1669_),
    .C1(_1670_),
    .D1(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__a22o_1 _5013_ (.A1(\mem[16][2] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][2] ),
    .X(_1673_));
 sky130_fd_sc_hd__a221o_1 _5014_ (.A1(\mem[6][2] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][2] ),
    .C1(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__a22o_1 _5015_ (.A1(\mem[28][2] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][2] ),
    .X(_1675_));
 sky130_fd_sc_hd__a221o_1 _5016_ (.A1(\mem[17][2] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][2] ),
    .C1(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__or4_4 _5017_ (.A(_1668_),
    .B(_1672_),
    .C(_1674_),
    .D(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_2 _5018_ (.A(_1677_),
    .X(net72));
 sky130_fd_sc_hd__and3_1 _5019_ (.A(_1589_),
    .B(\mem[24][3] ),
    .C(_1590_),
    .X(_1678_));
 sky130_fd_sc_hd__and3_1 _5020_ (.A(\mem[30][3] ),
    .B(_1543_),
    .C(_1592_),
    .X(_1679_));
 sky130_fd_sc_hd__and3_1 _5021_ (.A(_1594_),
    .B(\mem[27][3] ),
    .C(_1515_),
    .X(_1680_));
 sky130_fd_sc_hd__a2111o_1 _5022_ (.A1(\mem[12][3] ),
    .A2(_1512_),
    .B1(_1678_),
    .C1(_1679_),
    .D1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__and3_1 _5023_ (.A(_1599_),
    .B(\mem[15][3] ),
    .C(_1534_),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_4 _5024_ (.A(_1532_),
    .X(_1683_));
 sky130_fd_sc_hd__and3b_1 _5025_ (.A_N(_1601_),
    .B(_1683_),
    .C(\mem[13][3] ),
    .X(_1684_));
 sky130_fd_sc_hd__and3_1 _5026_ (.A(_1652_),
    .B(\mem[8][3] ),
    .C(_1523_),
    .X(_1685_));
 sky130_fd_sc_hd__a2111o_1 _5027_ (.A1(\mem[10][3] ),
    .A2(_1598_),
    .B1(_1682_),
    .C1(_1684_),
    .D1(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__inv_2 _5028_ (.A(\mem[3][3] ),
    .Y(_1687_));
 sky130_fd_sc_hd__buf_4 _5029_ (.A(_1549_),
    .X(_1688_));
 sky130_fd_sc_hd__nor3_1 _5030_ (.A(_1687_),
    .B(_1607_),
    .C(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__and4b_1 _5031_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][3] ),
    .D(_1610_),
    .X(_1690_));
 sky130_fd_sc_hd__and3b_1 _5032_ (.A_N(_1612_),
    .B(_1613_),
    .C(\mem[5][3] ),
    .X(_1691_));
 sky130_fd_sc_hd__a2111o_1 _5033_ (.A1(\mem[1][3] ),
    .A2(_1551_),
    .B1(_1689_),
    .C1(_1690_),
    .D1(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__and3_1 _5034_ (.A(\mem[18][3] ),
    .B(_1616_),
    .C(_1508_),
    .X(_1693_));
 sky130_fd_sc_hd__and3_1 _5035_ (.A(\mem[2][3] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1694_));
 sky130_fd_sc_hd__and3_1 _5036_ (.A(_1619_),
    .B(\mem[23][3] ),
    .C(_1573_),
    .X(_1695_));
 sky130_fd_sc_hd__a2111o_1 _5037_ (.A1(\mem[20][3] ),
    .A2(_1542_),
    .B1(_1693_),
    .C1(_1694_),
    .D1(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__or4_1 _5038_ (.A(_1681_),
    .B(_1686_),
    .C(_1692_),
    .D(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__a22o_1 _5039_ (.A1(\mem[7][3] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][3] ),
    .X(_1698_));
 sky130_fd_sc_hd__a22o_1 _5040_ (.A1(\mem[31][3] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][3] ),
    .X(_1699_));
 sky130_fd_sc_hd__a22o_1 _5041_ (.A1(\mem[11][3] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][3] ),
    .X(_1700_));
 sky130_fd_sc_hd__a2111o_1 _5042_ (.A1(\mem[26][3] ),
    .A2(_1624_),
    .B1(_1698_),
    .C1(_1699_),
    .D1(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__a22o_1 _5043_ (.A1(\mem[16][3] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][3] ),
    .X(_1702_));
 sky130_fd_sc_hd__a221o_1 _5044_ (.A1(\mem[6][3] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][3] ),
    .C1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__a22o_1 _5045_ (.A1(\mem[28][3] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][3] ),
    .X(_1704_));
 sky130_fd_sc_hd__a221o_1 _5046_ (.A1(\mem[17][3] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][3] ),
    .C1(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__or4_4 _5047_ (.A(_1697_),
    .B(_1701_),
    .C(_1703_),
    .D(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _5048_ (.A(_1706_),
    .X(net75));
 sky130_fd_sc_hd__and3_1 _5049_ (.A(_1589_),
    .B(\mem[24][4] ),
    .C(_1590_),
    .X(_1707_));
 sky130_fd_sc_hd__and3_1 _5050_ (.A(\mem[30][4] ),
    .B(_1543_),
    .C(_1592_),
    .X(_1708_));
 sky130_fd_sc_hd__and3_1 _5051_ (.A(_1594_),
    .B(\mem[27][4] ),
    .C(_1515_),
    .X(_1709_));
 sky130_fd_sc_hd__a2111o_1 _5052_ (.A1(\mem[12][4] ),
    .A2(_1512_),
    .B1(_1707_),
    .C1(_1708_),
    .D1(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__and3_1 _5053_ (.A(_1599_),
    .B(\mem[15][4] ),
    .C(_1534_),
    .X(_1711_));
 sky130_fd_sc_hd__and3b_1 _5054_ (.A_N(_1601_),
    .B(_1683_),
    .C(\mem[13][4] ),
    .X(_1712_));
 sky130_fd_sc_hd__and3_1 _5055_ (.A(_1652_),
    .B(\mem[8][4] ),
    .C(_1523_),
    .X(_1713_));
 sky130_fd_sc_hd__a2111o_1 _5056_ (.A1(\mem[10][4] ),
    .A2(_1598_),
    .B1(_1711_),
    .C1(_1712_),
    .D1(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__and4b_1 _5057_ (.A_N(_1655_),
    .B(_1656_),
    .C(\mem[22][4] ),
    .D(_1657_),
    .X(_1715_));
 sky130_fd_sc_hd__inv_2 _5058_ (.A(\mem[3][4] ),
    .Y(_1716_));
 sky130_fd_sc_hd__nor3_1 _5059_ (.A(_1716_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1717_));
 sky130_fd_sc_hd__buf_2 _5060_ (.A(_1532_),
    .X(_1718_));
 sky130_fd_sc_hd__and3b_1 _5061_ (.A_N(_1612_),
    .B(_1718_),
    .C(\mem[5][4] ),
    .X(_1719_));
 sky130_fd_sc_hd__a2111o_1 _5062_ (.A1(\mem[1][4] ),
    .A2(_1551_),
    .B1(_1715_),
    .C1(_1717_),
    .D1(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__and3_1 _5063_ (.A(\mem[18][4] ),
    .B(_1616_),
    .C(_1508_),
    .X(_1721_));
 sky130_fd_sc_hd__and3_1 _5064_ (.A(\mem[2][4] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1722_));
 sky130_fd_sc_hd__and3_1 _5065_ (.A(_1619_),
    .B(\mem[23][4] ),
    .C(_1573_),
    .X(_1723_));
 sky130_fd_sc_hd__a2111o_1 _5066_ (.A1(\mem[20][4] ),
    .A2(_1542_),
    .B1(_1721_),
    .C1(_1722_),
    .D1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__or4_1 _5067_ (.A(_1710_),
    .B(_1714_),
    .C(_1720_),
    .D(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__a22o_1 _5068_ (.A1(\mem[7][4] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][4] ),
    .X(_1726_));
 sky130_fd_sc_hd__a22o_1 _5069_ (.A1(\mem[31][4] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][4] ),
    .X(_1727_));
 sky130_fd_sc_hd__a22o_1 _5070_ (.A1(\mem[11][4] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][4] ),
    .X(_1728_));
 sky130_fd_sc_hd__a2111o_1 _5071_ (.A1(\mem[26][4] ),
    .A2(_1624_),
    .B1(_1726_),
    .C1(_1727_),
    .D1(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__a22o_1 _5072_ (.A1(\mem[16][4] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][4] ),
    .X(_1730_));
 sky130_fd_sc_hd__a221o_1 _5073_ (.A1(\mem[6][4] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][4] ),
    .C1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__a22o_1 _5074_ (.A1(\mem[28][4] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][4] ),
    .X(_1732_));
 sky130_fd_sc_hd__a221o_1 _5075_ (.A1(\mem[17][4] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][4] ),
    .C1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__or4_4 _5076_ (.A(_1725_),
    .B(_1729_),
    .C(_1731_),
    .D(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__buf_4 _5077_ (.A(_1734_),
    .X(net76));
 sky130_fd_sc_hd__and3_1 _5078_ (.A(_1589_),
    .B(\mem[24][5] ),
    .C(_1590_),
    .X(_1735_));
 sky130_fd_sc_hd__buf_4 _5079_ (.A(_1506_),
    .X(_1736_));
 sky130_fd_sc_hd__and3_1 _5080_ (.A(\mem[30][5] ),
    .B(_1543_),
    .C(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__and3_1 _5081_ (.A(_1594_),
    .B(\mem[27][5] ),
    .C(_1515_),
    .X(_1738_));
 sky130_fd_sc_hd__a2111o_1 _5082_ (.A1(\mem[12][5] ),
    .A2(_1512_),
    .B1(_1735_),
    .C1(_1737_),
    .D1(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_4 _5083_ (.A(_1532_),
    .X(_1740_));
 sky130_fd_sc_hd__and3_1 _5084_ (.A(_1740_),
    .B(\mem[15][5] ),
    .C(_1534_),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_4 _5085_ (.A(_1560_),
    .X(_1742_));
 sky130_fd_sc_hd__and3b_1 _5086_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][5] ),
    .X(_1743_));
 sky130_fd_sc_hd__and3_1 _5087_ (.A(_1652_),
    .B(\mem[8][5] ),
    .C(_1523_),
    .X(_1744_));
 sky130_fd_sc_hd__a2111o_1 _5088_ (.A1(\mem[10][5] ),
    .A2(_1598_),
    .B1(_1741_),
    .C1(_1743_),
    .D1(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__and4b_1 _5089_ (.A_N(_1655_),
    .B(_1656_),
    .C(\mem[22][5] ),
    .D(_1657_),
    .X(_1746_));
 sky130_fd_sc_hd__inv_2 _5090_ (.A(\mem[3][5] ),
    .Y(_1747_));
 sky130_fd_sc_hd__nor3_1 _5091_ (.A(_1747_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1748_));
 sky130_fd_sc_hd__buf_2 _5092_ (.A(_1556_),
    .X(_1749_));
 sky130_fd_sc_hd__and3b_1 _5093_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][5] ),
    .X(_1750_));
 sky130_fd_sc_hd__a2111o_1 _5094_ (.A1(\mem[1][5] ),
    .A2(_1551_),
    .B1(_1746_),
    .C1(_1748_),
    .D1(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__and3_1 _5095_ (.A(\mem[18][5] ),
    .B(_1616_),
    .C(_1508_),
    .X(_1752_));
 sky130_fd_sc_hd__and3_1 _5096_ (.A(\mem[2][5] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1753_));
 sky130_fd_sc_hd__and3_1 _5097_ (.A(_1619_),
    .B(\mem[23][5] ),
    .C(_1573_),
    .X(_1754_));
 sky130_fd_sc_hd__a2111o_1 _5098_ (.A1(\mem[20][5] ),
    .A2(_1542_),
    .B1(_1752_),
    .C1(_1753_),
    .D1(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__or4_1 _5099_ (.A(_1739_),
    .B(_1745_),
    .C(_1751_),
    .D(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__a22o_1 _5100_ (.A1(\mem[7][5] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][5] ),
    .X(_1757_));
 sky130_fd_sc_hd__a22o_1 _5101_ (.A1(\mem[31][5] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][5] ),
    .X(_1758_));
 sky130_fd_sc_hd__a22o_1 _5102_ (.A1(\mem[11][5] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][5] ),
    .X(_1759_));
 sky130_fd_sc_hd__a2111o_1 _5103_ (.A1(\mem[26][5] ),
    .A2(_1624_),
    .B1(_1757_),
    .C1(_1758_),
    .D1(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__a22o_1 _5104_ (.A1(\mem[16][5] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][5] ),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_1 _5105_ (.A1(\mem[6][5] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][5] ),
    .C1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__a22o_1 _5106_ (.A1(\mem[28][5] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][5] ),
    .X(_1763_));
 sky130_fd_sc_hd__a221o_1 _5107_ (.A1(\mem[17][5] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][5] ),
    .C1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__or4_4 _5108_ (.A(_1756_),
    .B(_1760_),
    .C(_1762_),
    .D(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__clkbuf_1 _5109_ (.A(_1765_),
    .X(net77));
 sky130_fd_sc_hd__and3_1 _5110_ (.A(_1589_),
    .B(\mem[24][6] ),
    .C(_1590_),
    .X(_1766_));
 sky130_fd_sc_hd__and3_1 _5111_ (.A(\mem[30][6] ),
    .B(_1543_),
    .C(_1736_),
    .X(_1767_));
 sky130_fd_sc_hd__and3_1 _5112_ (.A(_1594_),
    .B(\mem[27][6] ),
    .C(_1515_),
    .X(_1768_));
 sky130_fd_sc_hd__a2111o_1 _5113_ (.A1(\mem[12][6] ),
    .A2(_1512_),
    .B1(_1766_),
    .C1(_1767_),
    .D1(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__and3_1 _5114_ (.A(_1740_),
    .B(\mem[15][6] ),
    .C(_1534_),
    .X(_1770_));
 sky130_fd_sc_hd__and3b_1 _5115_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][6] ),
    .X(_1771_));
 sky130_fd_sc_hd__and3_1 _5116_ (.A(_1652_),
    .B(\mem[8][6] ),
    .C(_1523_),
    .X(_1772_));
 sky130_fd_sc_hd__a2111o_1 _5117_ (.A1(\mem[10][6] ),
    .A2(_1598_),
    .B1(_1770_),
    .C1(_1771_),
    .D1(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__and4b_1 _5118_ (.A_N(_1655_),
    .B(_1656_),
    .C(\mem[22][6] ),
    .D(_1657_),
    .X(_1774_));
 sky130_fd_sc_hd__inv_2 _5119_ (.A(\mem[3][6] ),
    .Y(_1775_));
 sky130_fd_sc_hd__nor3_1 _5120_ (.A(_1775_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1776_));
 sky130_fd_sc_hd__and3b_1 _5121_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][6] ),
    .X(_1777_));
 sky130_fd_sc_hd__a2111o_1 _5122_ (.A1(\mem[1][6] ),
    .A2(_1551_),
    .B1(_1774_),
    .C1(_1776_),
    .D1(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__clkbuf_4 _5123_ (.A(_1507_),
    .X(_1779_));
 sky130_fd_sc_hd__and3_1 _5124_ (.A(\mem[18][6] ),
    .B(_1616_),
    .C(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__and3_1 _5125_ (.A(\mem[2][6] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1781_));
 sky130_fd_sc_hd__and3_1 _5126_ (.A(_1619_),
    .B(\mem[23][6] ),
    .C(_1573_),
    .X(_1782_));
 sky130_fd_sc_hd__a2111o_1 _5127_ (.A1(\mem[20][6] ),
    .A2(_1542_),
    .B1(_1780_),
    .C1(_1781_),
    .D1(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__or4_1 _5128_ (.A(_1769_),
    .B(_1773_),
    .C(_1778_),
    .D(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__a22o_1 _5129_ (.A1(\mem[7][6] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][6] ),
    .X(_1785_));
 sky130_fd_sc_hd__a22o_1 _5130_ (.A1(\mem[31][6] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][6] ),
    .X(_1786_));
 sky130_fd_sc_hd__a22o_1 _5131_ (.A1(\mem[11][6] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][6] ),
    .X(_1787_));
 sky130_fd_sc_hd__a2111o_1 _5132_ (.A1(\mem[26][6] ),
    .A2(_1624_),
    .B1(_1785_),
    .C1(_1786_),
    .D1(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__a22o_1 _5133_ (.A1(\mem[16][6] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][6] ),
    .X(_1789_));
 sky130_fd_sc_hd__a221o_1 _5134_ (.A1(\mem[6][6] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][6] ),
    .C1(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__a22o_1 _5135_ (.A1(\mem[28][6] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][6] ),
    .X(_1791_));
 sky130_fd_sc_hd__a221o_1 _5136_ (.A1(\mem[17][6] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][6] ),
    .C1(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__or4_4 _5137_ (.A(_1784_),
    .B(_1788_),
    .C(_1790_),
    .D(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _5138_ (.A(_1793_),
    .X(net78));
 sky130_fd_sc_hd__and3_1 _5139_ (.A(_1589_),
    .B(\mem[24][7] ),
    .C(_1590_),
    .X(_1794_));
 sky130_fd_sc_hd__and3_1 _5140_ (.A(\mem[30][7] ),
    .B(_1543_),
    .C(_1736_),
    .X(_1795_));
 sky130_fd_sc_hd__and3_1 _5141_ (.A(_1594_),
    .B(\mem[27][7] ),
    .C(_1515_),
    .X(_1796_));
 sky130_fd_sc_hd__a2111o_1 _5142_ (.A1(\mem[12][7] ),
    .A2(_1512_),
    .B1(_1794_),
    .C1(_1795_),
    .D1(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__and3_1 _5143_ (.A(_1740_),
    .B(\mem[15][7] ),
    .C(_1534_),
    .X(_1798_));
 sky130_fd_sc_hd__and3b_1 _5144_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][7] ),
    .X(_1799_));
 sky130_fd_sc_hd__and3_1 _5145_ (.A(_1652_),
    .B(\mem[8][7] ),
    .C(_1523_),
    .X(_1800_));
 sky130_fd_sc_hd__a2111o_1 _5146_ (.A1(\mem[10][7] ),
    .A2(_1598_),
    .B1(_1798_),
    .C1(_1799_),
    .D1(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__inv_2 _5147_ (.A(\mem[3][7] ),
    .Y(_1802_));
 sky130_fd_sc_hd__nor3_1 _5148_ (.A(_1802_),
    .B(_1607_),
    .C(_1688_),
    .Y(_1803_));
 sky130_fd_sc_hd__and4b_1 _5149_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][7] ),
    .D(_1610_),
    .X(_1804_));
 sky130_fd_sc_hd__and3b_1 _5150_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][7] ),
    .X(_1805_));
 sky130_fd_sc_hd__a2111o_1 _5151_ (.A1(\mem[1][7] ),
    .A2(_1551_),
    .B1(_1803_),
    .C1(_1804_),
    .D1(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__clkbuf_4 _5152_ (.A(_1503_),
    .X(_1807_));
 sky130_fd_sc_hd__and3_1 _5153_ (.A(\mem[18][7] ),
    .B(_1807_),
    .C(_1779_),
    .X(_1808_));
 sky130_fd_sc_hd__and3_1 _5154_ (.A(\mem[2][7] ),
    .B(_1505_),
    .C(_1538_),
    .X(_1809_));
 sky130_fd_sc_hd__and3_1 _5155_ (.A(_1619_),
    .B(\mem[23][7] ),
    .C(_1573_),
    .X(_1810_));
 sky130_fd_sc_hd__a2111o_1 _5156_ (.A1(\mem[20][7] ),
    .A2(_1542_),
    .B1(_1808_),
    .C1(_1809_),
    .D1(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__or4_1 _5157_ (.A(_1797_),
    .B(_1801_),
    .C(_1806_),
    .D(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__a22o_1 _5158_ (.A1(\mem[7][7] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][7] ),
    .X(_1813_));
 sky130_fd_sc_hd__a22o_1 _5159_ (.A1(\mem[31][7] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][7] ),
    .X(_1814_));
 sky130_fd_sc_hd__a22o_1 _5160_ (.A1(\mem[11][7] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][7] ),
    .X(_1815_));
 sky130_fd_sc_hd__a2111o_1 _5161_ (.A1(\mem[26][7] ),
    .A2(_1624_),
    .B1(_1813_),
    .C1(_1814_),
    .D1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__a22o_1 _5162_ (.A1(\mem[16][7] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][7] ),
    .X(_1817_));
 sky130_fd_sc_hd__a221o_1 _5163_ (.A1(\mem[6][7] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][7] ),
    .C1(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__a22o_1 _5164_ (.A1(\mem[28][7] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][7] ),
    .X(_1819_));
 sky130_fd_sc_hd__a221o_1 _5165_ (.A1(\mem[17][7] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][7] ),
    .C1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__or4_1 _5166_ (.A(_1812_),
    .B(_1816_),
    .C(_1818_),
    .D(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__buf_4 _5167_ (.A(_1821_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 _5168_ (.A(_1519_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_4 _5169_ (.A(_1522_),
    .X(_1823_));
 sky130_fd_sc_hd__and3_1 _5170_ (.A(_1822_),
    .B(\mem[24][8] ),
    .C(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__and3_1 _5171_ (.A(\mem[30][8] ),
    .B(_1543_),
    .C(_1736_),
    .X(_1825_));
 sky130_fd_sc_hd__and3_1 _5172_ (.A(_1594_),
    .B(\mem[27][8] ),
    .C(_1515_),
    .X(_1826_));
 sky130_fd_sc_hd__a2111o_1 _5173_ (.A1(\mem[12][8] ),
    .A2(_1512_),
    .B1(_1824_),
    .C1(_1825_),
    .D1(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__and3_1 _5174_ (.A(_1740_),
    .B(\mem[15][8] ),
    .C(_1534_),
    .X(_1828_));
 sky130_fd_sc_hd__and3b_1 _5175_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][8] ),
    .X(_1829_));
 sky130_fd_sc_hd__and3_1 _5176_ (.A(_1652_),
    .B(\mem[8][8] ),
    .C(_1523_),
    .X(_1830_));
 sky130_fd_sc_hd__a2111o_1 _5177_ (.A1(\mem[10][8] ),
    .A2(_1598_),
    .B1(_1828_),
    .C1(_1829_),
    .D1(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__and4b_1 _5178_ (.A_N(_1655_),
    .B(_1656_),
    .C(\mem[22][8] ),
    .D(_1507_),
    .X(_1832_));
 sky130_fd_sc_hd__inv_2 _5179_ (.A(\mem[3][8] ),
    .Y(_1833_));
 sky130_fd_sc_hd__nor3_1 _5180_ (.A(_1833_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1834_));
 sky130_fd_sc_hd__and3b_1 _5181_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][8] ),
    .X(_1835_));
 sky130_fd_sc_hd__a2111o_1 _5182_ (.A1(\mem[1][8] ),
    .A2(_1551_),
    .B1(_1832_),
    .C1(_1834_),
    .D1(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__and3_1 _5183_ (.A(\mem[18][8] ),
    .B(_1807_),
    .C(_1779_),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_4 _5184_ (.A(_1504_),
    .X(_1838_));
 sky130_fd_sc_hd__buf_4 _5185_ (.A(_1524_),
    .X(_1839_));
 sky130_fd_sc_hd__and3_1 _5186_ (.A(\mem[2][8] ),
    .B(_1838_),
    .C(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__and3_1 _5187_ (.A(_1619_),
    .B(\mem[23][8] ),
    .C(_1573_),
    .X(_1841_));
 sky130_fd_sc_hd__a2111o_1 _5188_ (.A1(\mem[20][8] ),
    .A2(_1542_),
    .B1(_1837_),
    .C1(_1840_),
    .D1(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__or4_1 _5189_ (.A(_1827_),
    .B(_1831_),
    .C(_1836_),
    .D(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__a22o_1 _5190_ (.A1(\mem[7][8] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][8] ),
    .X(_1844_));
 sky130_fd_sc_hd__a22o_1 _5191_ (.A1(\mem[31][8] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][8] ),
    .X(_1845_));
 sky130_fd_sc_hd__a22o_1 _5192_ (.A1(\mem[11][8] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][8] ),
    .X(_1846_));
 sky130_fd_sc_hd__a2111o_1 _5193_ (.A1(\mem[26][8] ),
    .A2(_1624_),
    .B1(_1844_),
    .C1(_1845_),
    .D1(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__a22o_1 _5194_ (.A1(\mem[16][8] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][8] ),
    .X(_1848_));
 sky130_fd_sc_hd__a221o_1 _5195_ (.A1(\mem[6][8] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][8] ),
    .C1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__a22o_1 _5196_ (.A1(\mem[28][8] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][8] ),
    .X(_1850_));
 sky130_fd_sc_hd__a221o_1 _5197_ (.A1(\mem[17][8] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][8] ),
    .C1(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__or4_4 _5198_ (.A(_1843_),
    .B(_1847_),
    .C(_1849_),
    .D(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_1 _5199_ (.A(_1852_),
    .X(net80));
 sky130_fd_sc_hd__and3_1 _5200_ (.A(_1822_),
    .B(\mem[24][9] ),
    .C(_1823_),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_4 _5201_ (.A(_1509_),
    .X(_1854_));
 sky130_fd_sc_hd__and3_1 _5202_ (.A(\mem[30][9] ),
    .B(_1854_),
    .C(_1736_),
    .X(_1855_));
 sky130_fd_sc_hd__clkbuf_4 _5203_ (.A(_1519_),
    .X(_1856_));
 sky130_fd_sc_hd__and3_1 _5204_ (.A(_1856_),
    .B(\mem[27][9] ),
    .C(_1515_),
    .X(_1857_));
 sky130_fd_sc_hd__a2111o_1 _5205_ (.A1(\mem[12][9] ),
    .A2(_1512_),
    .B1(_1853_),
    .C1(_1855_),
    .D1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__and3_1 _5206_ (.A(_1740_),
    .B(\mem[15][9] ),
    .C(_1534_),
    .X(_1859_));
 sky130_fd_sc_hd__and3b_1 _5207_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][9] ),
    .X(_1860_));
 sky130_fd_sc_hd__clkbuf_4 _5208_ (.A(_1522_),
    .X(_1861_));
 sky130_fd_sc_hd__and3_1 _5209_ (.A(_1652_),
    .B(\mem[8][9] ),
    .C(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__a2111o_1 _5210_ (.A1(\mem[10][9] ),
    .A2(_1598_),
    .B1(_1859_),
    .C1(_1860_),
    .D1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__inv_2 _5211_ (.A(\mem[3][9] ),
    .Y(_1864_));
 sky130_fd_sc_hd__nor3_1 _5212_ (.A(_1864_),
    .B(_1607_),
    .C(_1688_),
    .Y(_1865_));
 sky130_fd_sc_hd__and4b_1 _5213_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][9] ),
    .D(_1610_),
    .X(_1866_));
 sky130_fd_sc_hd__and3b_1 _5214_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][9] ),
    .X(_1867_));
 sky130_fd_sc_hd__a2111o_1 _5215_ (.A1(\mem[1][9] ),
    .A2(_1551_),
    .B1(_1865_),
    .C1(_1866_),
    .D1(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__and3_1 _5216_ (.A(\mem[18][9] ),
    .B(_1807_),
    .C(_1779_),
    .X(_1869_));
 sky130_fd_sc_hd__and3_1 _5217_ (.A(\mem[2][9] ),
    .B(_1838_),
    .C(_1839_),
    .X(_1870_));
 sky130_fd_sc_hd__and3_1 _5218_ (.A(_1619_),
    .B(\mem[23][9] ),
    .C(_1573_),
    .X(_1871_));
 sky130_fd_sc_hd__a2111o_1 _5219_ (.A1(\mem[20][9] ),
    .A2(_1542_),
    .B1(_1869_),
    .C1(_1870_),
    .D1(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__or4_1 _5220_ (.A(_1858_),
    .B(_1863_),
    .C(_1868_),
    .D(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__a22o_1 _5221_ (.A1(\mem[7][9] ),
    .A2(_1566_),
    .B1(_1572_),
    .B2(\mem[9][9] ),
    .X(_1874_));
 sky130_fd_sc_hd__a22o_1 _5222_ (.A1(\mem[31][9] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][9] ),
    .X(_1875_));
 sky130_fd_sc_hd__a22o_1 _5223_ (.A1(\mem[11][9] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][9] ),
    .X(_1876_));
 sky130_fd_sc_hd__a2111o_1 _5224_ (.A1(\mem[26][9] ),
    .A2(_1624_),
    .B1(_1874_),
    .C1(_1875_),
    .D1(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__a22o_1 _5225_ (.A1(\mem[16][9] ),
    .A2(_1547_),
    .B1(_1581_),
    .B2(\mem[19][9] ),
    .X(_1878_));
 sky130_fd_sc_hd__a221o_1 _5226_ (.A1(\mem[6][9] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][9] ),
    .C1(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__a22o_1 _5227_ (.A1(\mem[28][9] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][9] ),
    .X(_1880_));
 sky130_fd_sc_hd__a221o_1 _5228_ (.A1(\mem[17][9] ),
    .A2(_1531_),
    .B1(_1638_),
    .B2(\mem[21][9] ),
    .C1(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__or4_4 _5229_ (.A(_1873_),
    .B(_1877_),
    .C(_1879_),
    .D(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__clkbuf_1 _5230_ (.A(_1882_),
    .X(net81));
 sky130_fd_sc_hd__buf_4 _5231_ (.A(_1511_),
    .X(_1883_));
 sky130_fd_sc_hd__and3_1 _5232_ (.A(_1822_),
    .B(\mem[24][10] ),
    .C(_1823_),
    .X(_1884_));
 sky130_fd_sc_hd__and3_1 _5233_ (.A(\mem[30][10] ),
    .B(_1854_),
    .C(_1736_),
    .X(_1885_));
 sky130_fd_sc_hd__clkbuf_4 _5234_ (.A(_1497_),
    .X(_1886_));
 sky130_fd_sc_hd__and3_1 _5235_ (.A(_1856_),
    .B(\mem[27][10] ),
    .C(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__a2111o_1 _5236_ (.A1(\mem[12][10] ),
    .A2(_1883_),
    .B1(_1884_),
    .C1(_1885_),
    .D1(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__clkbuf_4 _5237_ (.A(_1500_),
    .X(_1889_));
 sky130_fd_sc_hd__and3_1 _5238_ (.A(_1740_),
    .B(\mem[15][10] ),
    .C(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__and3b_1 _5239_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][10] ),
    .X(_1891_));
 sky130_fd_sc_hd__and3_1 _5240_ (.A(_1652_),
    .B(\mem[8][10] ),
    .C(_1861_),
    .X(_1892_));
 sky130_fd_sc_hd__a2111o_1 _5241_ (.A1(\mem[10][10] ),
    .A2(_1598_),
    .B1(_1890_),
    .C1(_1891_),
    .D1(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__buf_4 _5242_ (.A(_1550_),
    .X(_1894_));
 sky130_fd_sc_hd__and4b_1 _5243_ (.A_N(_1655_),
    .B(_1656_),
    .C(\mem[22][10] ),
    .D(_1507_),
    .X(_1895_));
 sky130_fd_sc_hd__inv_2 _5244_ (.A(\mem[3][10] ),
    .Y(_1896_));
 sky130_fd_sc_hd__nor3_1 _5245_ (.A(_1896_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1897_));
 sky130_fd_sc_hd__and3b_1 _5246_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][10] ),
    .X(_1898_));
 sky130_fd_sc_hd__a2111o_1 _5247_ (.A1(\mem[1][10] ),
    .A2(_1894_),
    .B1(_1895_),
    .C1(_1897_),
    .D1(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__buf_4 _5248_ (.A(_1541_),
    .X(_1900_));
 sky130_fd_sc_hd__and3_1 _5249_ (.A(\mem[18][10] ),
    .B(_1807_),
    .C(_1779_),
    .X(_1901_));
 sky130_fd_sc_hd__and3_1 _5250_ (.A(\mem[2][10] ),
    .B(_1838_),
    .C(_1839_),
    .X(_1902_));
 sky130_fd_sc_hd__clkbuf_4 _5251_ (.A(_1519_),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_4 _5252_ (.A(_1564_),
    .X(_1904_));
 sky130_fd_sc_hd__and3_1 _5253_ (.A(_1903_),
    .B(\mem[23][10] ),
    .C(_1904_),
    .X(_1905_));
 sky130_fd_sc_hd__a2111o_1 _5254_ (.A1(\mem[20][10] ),
    .A2(_1900_),
    .B1(_1901_),
    .C1(_1902_),
    .D1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__or4_1 _5255_ (.A(_1888_),
    .B(_1893_),
    .C(_1899_),
    .D(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_8 _5256_ (.A(_1565_),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_8 _5257_ (.A(_1571_),
    .X(_1909_));
 sky130_fd_sc_hd__a22o_1 _5258_ (.A1(\mem[7][10] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][10] ),
    .X(_1910_));
 sky130_fd_sc_hd__a22o_1 _5259_ (.A1(\mem[31][10] ),
    .A2(_1626_),
    .B1(_1627_),
    .B2(\mem[25][10] ),
    .X(_1911_));
 sky130_fd_sc_hd__a22o_1 _5260_ (.A1(\mem[11][10] ),
    .A2(_1629_),
    .B1(_1630_),
    .B2(\mem[14][10] ),
    .X(_1912_));
 sky130_fd_sc_hd__a2111o_1 _5261_ (.A1(\mem[26][10] ),
    .A2(_1624_),
    .B1(_1910_),
    .C1(_1911_),
    .D1(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__buf_6 _5262_ (.A(_1546_),
    .X(_1914_));
 sky130_fd_sc_hd__buf_6 _5263_ (.A(_1580_),
    .X(_1915_));
 sky130_fd_sc_hd__a22o_1 _5264_ (.A1(\mem[16][10] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][10] ),
    .X(_1916_));
 sky130_fd_sc_hd__a221o_1 _5265_ (.A1(\mem[6][10] ),
    .A2(_1633_),
    .B1(_1634_),
    .B2(\mem[4][10] ),
    .C1(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__buf_6 _5266_ (.A(_1530_),
    .X(_1918_));
 sky130_fd_sc_hd__a22o_1 _5267_ (.A1(\mem[28][10] ),
    .A2(_1640_),
    .B1(_1642_),
    .B2(\mem[29][10] ),
    .X(_1919_));
 sky130_fd_sc_hd__a221o_1 _5268_ (.A1(\mem[17][10] ),
    .A2(_1918_),
    .B1(_1638_),
    .B2(\mem[21][10] ),
    .C1(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__or4_2 _5269_ (.A(_1907_),
    .B(_1913_),
    .C(_1917_),
    .D(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__buf_4 _5270_ (.A(_1921_),
    .X(net51));
 sky130_fd_sc_hd__and3_1 _5271_ (.A(_1822_),
    .B(\mem[24][11] ),
    .C(_1823_),
    .X(_1922_));
 sky130_fd_sc_hd__and3_1 _5272_ (.A(\mem[30][11] ),
    .B(_1854_),
    .C(_1736_),
    .X(_1923_));
 sky130_fd_sc_hd__and3_1 _5273_ (.A(_1856_),
    .B(\mem[27][11] ),
    .C(_1886_),
    .X(_1924_));
 sky130_fd_sc_hd__a2111o_1 _5274_ (.A1(\mem[12][11] ),
    .A2(_1883_),
    .B1(_1922_),
    .C1(_1923_),
    .D1(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__buf_4 _5275_ (.A(_1597_),
    .X(_1926_));
 sky130_fd_sc_hd__and3_1 _5276_ (.A(_1740_),
    .B(\mem[15][11] ),
    .C(_1889_),
    .X(_1927_));
 sky130_fd_sc_hd__and3b_1 _5277_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][11] ),
    .X(_1928_));
 sky130_fd_sc_hd__and3_1 _5278_ (.A(_1652_),
    .B(\mem[8][11] ),
    .C(_1861_),
    .X(_1929_));
 sky130_fd_sc_hd__a2111o_1 _5279_ (.A1(\mem[10][11] ),
    .A2(_1926_),
    .B1(_1927_),
    .C1(_1928_),
    .D1(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__clkbuf_4 _5280_ (.A(_1517_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_4 _5281_ (.A(_1516_),
    .X(_1932_));
 sky130_fd_sc_hd__and4b_1 _5282_ (.A_N(_1931_),
    .B(_1932_),
    .C(\mem[22][11] ),
    .D(_1507_),
    .X(_1933_));
 sky130_fd_sc_hd__inv_2 _5283_ (.A(\mem[3][11] ),
    .Y(_1934_));
 sky130_fd_sc_hd__nor3_1 _5284_ (.A(_1934_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1935_));
 sky130_fd_sc_hd__and3b_1 _5285_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][11] ),
    .X(_1936_));
 sky130_fd_sc_hd__a2111o_1 _5286_ (.A1(\mem[1][11] ),
    .A2(_1894_),
    .B1(_1933_),
    .C1(_1935_),
    .D1(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__and3_1 _5287_ (.A(\mem[18][11] ),
    .B(_1807_),
    .C(_1779_),
    .X(_1938_));
 sky130_fd_sc_hd__and3_1 _5288_ (.A(\mem[2][11] ),
    .B(_1838_),
    .C(_1839_),
    .X(_1939_));
 sky130_fd_sc_hd__and3_1 _5289_ (.A(_1903_),
    .B(\mem[23][11] ),
    .C(_1904_),
    .X(_1940_));
 sky130_fd_sc_hd__a2111o_1 _5290_ (.A1(\mem[20][11] ),
    .A2(_1900_),
    .B1(_1938_),
    .C1(_1939_),
    .D1(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__or4_1 _5291_ (.A(_1925_),
    .B(_1930_),
    .C(_1937_),
    .D(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__buf_6 _5292_ (.A(_1623_),
    .X(_1943_));
 sky130_fd_sc_hd__a22o_1 _5293_ (.A1(\mem[7][11] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][11] ),
    .X(_1944_));
 sky130_fd_sc_hd__buf_6 _5294_ (.A(_1501_),
    .X(_1945_));
 sky130_fd_sc_hd__buf_6 _5295_ (.A(_1520_),
    .X(_1946_));
 sky130_fd_sc_hd__a22o_1 _5296_ (.A1(\mem[31][11] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][11] ),
    .X(_1947_));
 sky130_fd_sc_hd__buf_6 _5297_ (.A(_1498_),
    .X(_1948_));
 sky130_fd_sc_hd__buf_6 _5298_ (.A(_1525_),
    .X(_1949_));
 sky130_fd_sc_hd__a22o_1 _5299_ (.A1(\mem[11][11] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][11] ),
    .X(_1950_));
 sky130_fd_sc_hd__a2111o_1 _5300_ (.A1(\mem[26][11] ),
    .A2(_1943_),
    .B1(_1944_),
    .C1(_1947_),
    .D1(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__buf_6 _5301_ (.A(_1539_),
    .X(_1952_));
 sky130_fd_sc_hd__buf_6 _5302_ (.A(_1554_),
    .X(_1953_));
 sky130_fd_sc_hd__a22o_1 _5303_ (.A1(\mem[16][11] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][11] ),
    .X(_1954_));
 sky130_fd_sc_hd__a221o_1 _5304_ (.A1(\mem[6][11] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][11] ),
    .C1(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__buf_6 _5305_ (.A(_1637_),
    .X(_1956_));
 sky130_fd_sc_hd__buf_6 _5306_ (.A(_1639_),
    .X(_1957_));
 sky130_fd_sc_hd__buf_6 _5307_ (.A(_1641_),
    .X(_1958_));
 sky130_fd_sc_hd__a22o_1 _5308_ (.A1(\mem[28][11] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][11] ),
    .X(_1959_));
 sky130_fd_sc_hd__a221o_1 _5309_ (.A1(\mem[17][11] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][11] ),
    .C1(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__or4_4 _5310_ (.A(_1942_),
    .B(_1951_),
    .C(_1955_),
    .D(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__clkbuf_1 _5311_ (.A(_1961_),
    .X(net52));
 sky130_fd_sc_hd__and3_1 _5312_ (.A(_1822_),
    .B(\mem[24][12] ),
    .C(_1823_),
    .X(_1962_));
 sky130_fd_sc_hd__and3_1 _5313_ (.A(\mem[30][12] ),
    .B(_1854_),
    .C(_1736_),
    .X(_1963_));
 sky130_fd_sc_hd__and3_1 _5314_ (.A(_1856_),
    .B(\mem[27][12] ),
    .C(_1886_),
    .X(_1964_));
 sky130_fd_sc_hd__a2111o_1 _5315_ (.A1(\mem[12][12] ),
    .A2(_1883_),
    .B1(_1962_),
    .C1(_1963_),
    .D1(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__and3_1 _5316_ (.A(_1740_),
    .B(\mem[15][12] ),
    .C(_1889_),
    .X(_1966_));
 sky130_fd_sc_hd__and3b_1 _5317_ (.A_N(_1742_),
    .B(_1683_),
    .C(\mem[13][12] ),
    .X(_1967_));
 sky130_fd_sc_hd__and3_1 _5318_ (.A(_1613_),
    .B(\mem[8][12] ),
    .C(_1861_),
    .X(_1968_));
 sky130_fd_sc_hd__a2111o_1 _5319_ (.A1(\mem[10][12] ),
    .A2(_1926_),
    .B1(_1966_),
    .C1(_1967_),
    .D1(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__and4b_1 _5320_ (.A_N(_1931_),
    .B(_1932_),
    .C(\mem[22][12] ),
    .D(_1507_),
    .X(_1970_));
 sky130_fd_sc_hd__inv_2 _5321_ (.A(\mem[3][12] ),
    .Y(_1971_));
 sky130_fd_sc_hd__nor3_1 _5322_ (.A(_1971_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1972_));
 sky130_fd_sc_hd__and3b_1 _5323_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][12] ),
    .X(_1973_));
 sky130_fd_sc_hd__a2111o_1 _5324_ (.A1(\mem[1][12] ),
    .A2(_1894_),
    .B1(_1970_),
    .C1(_1972_),
    .D1(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__and3_1 _5325_ (.A(\mem[18][12] ),
    .B(_1807_),
    .C(_1779_),
    .X(_1975_));
 sky130_fd_sc_hd__and3_1 _5326_ (.A(\mem[2][12] ),
    .B(_1838_),
    .C(_1839_),
    .X(_1976_));
 sky130_fd_sc_hd__and3_1 _5327_ (.A(_1903_),
    .B(\mem[23][12] ),
    .C(_1904_),
    .X(_1977_));
 sky130_fd_sc_hd__a2111o_1 _5328_ (.A1(\mem[20][12] ),
    .A2(_1900_),
    .B1(_1975_),
    .C1(_1976_),
    .D1(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__or4_1 _5329_ (.A(_1965_),
    .B(_1969_),
    .C(_1974_),
    .D(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__a22o_1 _5330_ (.A1(\mem[7][12] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][12] ),
    .X(_1980_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(\mem[31][12] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][12] ),
    .X(_1981_));
 sky130_fd_sc_hd__a22o_1 _5332_ (.A1(\mem[11][12] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][12] ),
    .X(_1982_));
 sky130_fd_sc_hd__a2111o_1 _5333_ (.A1(\mem[26][12] ),
    .A2(_1943_),
    .B1(_1980_),
    .C1(_1981_),
    .D1(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__a22o_1 _5334_ (.A1(\mem[16][12] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][12] ),
    .X(_1984_));
 sky130_fd_sc_hd__a221o_1 _5335_ (.A1(\mem[6][12] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][12] ),
    .C1(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__a22o_1 _5336_ (.A1(\mem[28][12] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][12] ),
    .X(_1986_));
 sky130_fd_sc_hd__a221o_1 _5337_ (.A1(\mem[17][12] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][12] ),
    .C1(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__or4_4 _5338_ (.A(_1979_),
    .B(_1983_),
    .C(_1985_),
    .D(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__clkbuf_2 _5339_ (.A(_1988_),
    .X(net53));
 sky130_fd_sc_hd__and3_1 _5340_ (.A(_1822_),
    .B(\mem[24][13] ),
    .C(_1823_),
    .X(_1989_));
 sky130_fd_sc_hd__and3_1 _5341_ (.A(\mem[30][13] ),
    .B(_1854_),
    .C(_1736_),
    .X(_1990_));
 sky130_fd_sc_hd__and3_1 _5342_ (.A(_1856_),
    .B(\mem[27][13] ),
    .C(_1886_),
    .X(_1991_));
 sky130_fd_sc_hd__a2111o_1 _5343_ (.A1(\mem[12][13] ),
    .A2(_1883_),
    .B1(_1989_),
    .C1(_1990_),
    .D1(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__and3_1 _5344_ (.A(_1740_),
    .B(\mem[15][13] ),
    .C(_1889_),
    .X(_1993_));
 sky130_fd_sc_hd__and3b_1 _5345_ (.A_N(_1742_),
    .B(_1599_),
    .C(\mem[13][13] ),
    .X(_1994_));
 sky130_fd_sc_hd__and3_1 _5346_ (.A(_1613_),
    .B(\mem[8][13] ),
    .C(_1861_),
    .X(_1995_));
 sky130_fd_sc_hd__a2111o_1 _5347_ (.A1(\mem[10][13] ),
    .A2(_1926_),
    .B1(_1993_),
    .C1(_1994_),
    .D1(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__and4b_1 _5348_ (.A_N(_1931_),
    .B(_1932_),
    .C(\mem[22][13] ),
    .D(_1507_),
    .X(_1997_));
 sky130_fd_sc_hd__inv_2 _5349_ (.A(\mem[3][13] ),
    .Y(_1998_));
 sky130_fd_sc_hd__nor3_1 _5350_ (.A(_1998_),
    .B(_1584_),
    .C(_1660_),
    .Y(_1999_));
 sky130_fd_sc_hd__and3b_1 _5351_ (.A_N(_1749_),
    .B(_1718_),
    .C(\mem[5][13] ),
    .X(_2000_));
 sky130_fd_sc_hd__a2111o_1 _5352_ (.A1(\mem[1][13] ),
    .A2(_1894_),
    .B1(_1997_),
    .C1(_1999_),
    .D1(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__and3_1 _5353_ (.A(\mem[18][13] ),
    .B(_1807_),
    .C(_1779_),
    .X(_2002_));
 sky130_fd_sc_hd__and3_1 _5354_ (.A(\mem[2][13] ),
    .B(_1838_),
    .C(_1839_),
    .X(_2003_));
 sky130_fd_sc_hd__and3_1 _5355_ (.A(_1903_),
    .B(\mem[23][13] ),
    .C(_1904_),
    .X(_2004_));
 sky130_fd_sc_hd__a2111o_1 _5356_ (.A1(\mem[20][13] ),
    .A2(_1900_),
    .B1(_2002_),
    .C1(_2003_),
    .D1(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__or4_1 _5357_ (.A(_1992_),
    .B(_1996_),
    .C(_2001_),
    .D(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__a22o_1 _5358_ (.A1(\mem[7][13] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][13] ),
    .X(_2007_));
 sky130_fd_sc_hd__a22o_1 _5359_ (.A1(\mem[31][13] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][13] ),
    .X(_2008_));
 sky130_fd_sc_hd__a22o_1 _5360_ (.A1(\mem[11][13] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][13] ),
    .X(_2009_));
 sky130_fd_sc_hd__a2111o_1 _5361_ (.A1(\mem[26][13] ),
    .A2(_1943_),
    .B1(_2007_),
    .C1(_2008_),
    .D1(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__a22o_1 _5362_ (.A1(\mem[16][13] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][13] ),
    .X(_2011_));
 sky130_fd_sc_hd__a221o_1 _5363_ (.A1(\mem[6][13] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][13] ),
    .C1(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__a22o_1 _5364_ (.A1(\mem[28][13] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][13] ),
    .X(_2013_));
 sky130_fd_sc_hd__a221o_1 _5365_ (.A1(\mem[17][13] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][13] ),
    .C1(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__or4_4 _5366_ (.A(_2006_),
    .B(_2010_),
    .C(_2012_),
    .D(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__clkbuf_1 _5367_ (.A(_2015_),
    .X(net54));
 sky130_fd_sc_hd__and3_1 _5368_ (.A(_1822_),
    .B(\mem[24][14] ),
    .C(_1823_),
    .X(_2016_));
 sky130_fd_sc_hd__and3_1 _5369_ (.A(\mem[30][14] ),
    .B(_1854_),
    .C(_1736_),
    .X(_2017_));
 sky130_fd_sc_hd__and3_1 _5370_ (.A(_1856_),
    .B(\mem[27][14] ),
    .C(_1886_),
    .X(_2018_));
 sky130_fd_sc_hd__a2111o_1 _5371_ (.A1(\mem[12][14] ),
    .A2(_1883_),
    .B1(_2016_),
    .C1(_2017_),
    .D1(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__and3_1 _5372_ (.A(_1740_),
    .B(\mem[15][14] ),
    .C(_1889_),
    .X(_2020_));
 sky130_fd_sc_hd__and3b_1 _5373_ (.A_N(_1742_),
    .B(_1599_),
    .C(\mem[13][14] ),
    .X(_2021_));
 sky130_fd_sc_hd__and3_1 _5374_ (.A(_1613_),
    .B(\mem[8][14] ),
    .C(_1861_),
    .X(_2022_));
 sky130_fd_sc_hd__a2111o_1 _5375_ (.A1(\mem[10][14] ),
    .A2(_1926_),
    .B1(_2020_),
    .C1(_2021_),
    .D1(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__and4b_1 _5376_ (.A_N(_1931_),
    .B(_1932_),
    .C(\mem[22][14] ),
    .D(_1507_),
    .X(_2024_));
 sky130_fd_sc_hd__inv_2 _5377_ (.A(\mem[3][14] ),
    .Y(_2025_));
 sky130_fd_sc_hd__buf_4 _5378_ (.A(_1579_),
    .X(_2026_));
 sky130_fd_sc_hd__nor3_1 _5379_ (.A(_2025_),
    .B(_2026_),
    .C(_1660_),
    .Y(_2027_));
 sky130_fd_sc_hd__clkbuf_4 _5380_ (.A(_1532_),
    .X(_2028_));
 sky130_fd_sc_hd__and3b_1 _5381_ (.A_N(_1749_),
    .B(_2028_),
    .C(\mem[5][14] ),
    .X(_2029_));
 sky130_fd_sc_hd__a2111o_1 _5382_ (.A1(\mem[1][14] ),
    .A2(_1894_),
    .B1(_2024_),
    .C1(_2027_),
    .D1(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__and3_1 _5383_ (.A(\mem[18][14] ),
    .B(_1807_),
    .C(_1779_),
    .X(_2031_));
 sky130_fd_sc_hd__and3_1 _5384_ (.A(\mem[2][14] ),
    .B(_1838_),
    .C(_1839_),
    .X(_2032_));
 sky130_fd_sc_hd__and3_1 _5385_ (.A(_1903_),
    .B(\mem[23][14] ),
    .C(_1904_),
    .X(_2033_));
 sky130_fd_sc_hd__a2111o_1 _5386_ (.A1(\mem[20][14] ),
    .A2(_1900_),
    .B1(_2031_),
    .C1(_2032_),
    .D1(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__or4_1 _5387_ (.A(_2019_),
    .B(_2023_),
    .C(_2030_),
    .D(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__a22o_1 _5388_ (.A1(\mem[7][14] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][14] ),
    .X(_2036_));
 sky130_fd_sc_hd__a22o_1 _5389_ (.A1(\mem[31][14] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][14] ),
    .X(_2037_));
 sky130_fd_sc_hd__a22o_1 _5390_ (.A1(\mem[11][14] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][14] ),
    .X(_2038_));
 sky130_fd_sc_hd__a2111o_1 _5391_ (.A1(\mem[26][14] ),
    .A2(_1943_),
    .B1(_2036_),
    .C1(_2037_),
    .D1(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__a22o_1 _5392_ (.A1(\mem[16][14] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][14] ),
    .X(_2040_));
 sky130_fd_sc_hd__a221o_1 _5393_ (.A1(\mem[6][14] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][14] ),
    .C1(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__a22o_1 _5394_ (.A1(\mem[28][14] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][14] ),
    .X(_2042_));
 sky130_fd_sc_hd__a221o_1 _5395_ (.A1(\mem[17][14] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][14] ),
    .C1(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__or4_4 _5396_ (.A(_2035_),
    .B(_2039_),
    .C(_2041_),
    .D(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _5397_ (.A(_2044_),
    .X(net55));
 sky130_fd_sc_hd__and3_1 _5398_ (.A(_1822_),
    .B(\mem[24][15] ),
    .C(_1823_),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_4 _5399_ (.A(_1506_),
    .X(_2046_));
 sky130_fd_sc_hd__and3_1 _5400_ (.A(\mem[30][15] ),
    .B(_1854_),
    .C(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__and3_1 _5401_ (.A(_1856_),
    .B(\mem[27][15] ),
    .C(_1886_),
    .X(_2048_));
 sky130_fd_sc_hd__a2111o_1 _5402_ (.A1(\mem[12][15] ),
    .A2(_1883_),
    .B1(_2045_),
    .C1(_2047_),
    .D1(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_4 _5403_ (.A(_1493_),
    .X(_2050_));
 sky130_fd_sc_hd__and3_1 _5404_ (.A(_2050_),
    .B(\mem[15][15] ),
    .C(_1889_),
    .X(_2051_));
 sky130_fd_sc_hd__and3b_1 _5405_ (.A_N(_1560_),
    .B(_1599_),
    .C(\mem[13][15] ),
    .X(_2052_));
 sky130_fd_sc_hd__and3_1 _5406_ (.A(_1613_),
    .B(\mem[8][15] ),
    .C(_1861_),
    .X(_2053_));
 sky130_fd_sc_hd__a2111o_1 _5407_ (.A1(\mem[10][15] ),
    .A2(_1926_),
    .B1(_2051_),
    .C1(_2052_),
    .D1(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__and4b_1 _5408_ (.A_N(_1931_),
    .B(_1932_),
    .C(\mem[22][15] ),
    .D(_1507_),
    .X(_2055_));
 sky130_fd_sc_hd__inv_2 _5409_ (.A(\mem[3][15] ),
    .Y(_2056_));
 sky130_fd_sc_hd__nor3_1 _5410_ (.A(_2056_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2057_));
 sky130_fd_sc_hd__and3b_1 _5411_ (.A_N(_1556_),
    .B(_2028_),
    .C(\mem[5][15] ),
    .X(_2058_));
 sky130_fd_sc_hd__a2111o_1 _5412_ (.A1(\mem[1][15] ),
    .A2(_1894_),
    .B1(_2055_),
    .C1(_2057_),
    .D1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__and3_1 _5413_ (.A(\mem[18][15] ),
    .B(_1807_),
    .C(_1779_),
    .X(_2060_));
 sky130_fd_sc_hd__and3_1 _5414_ (.A(\mem[2][15] ),
    .B(_1838_),
    .C(_1839_),
    .X(_2061_));
 sky130_fd_sc_hd__and3_1 _5415_ (.A(_1903_),
    .B(\mem[23][15] ),
    .C(_1904_),
    .X(_2062_));
 sky130_fd_sc_hd__a2111o_1 _5416_ (.A1(\mem[20][15] ),
    .A2(_1900_),
    .B1(_2060_),
    .C1(_2061_),
    .D1(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__or4_1 _5417_ (.A(_2049_),
    .B(_2054_),
    .C(_2059_),
    .D(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__a22o_1 _5418_ (.A1(\mem[7][15] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][15] ),
    .X(_2065_));
 sky130_fd_sc_hd__a22o_1 _5419_ (.A1(\mem[31][15] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][15] ),
    .X(_2066_));
 sky130_fd_sc_hd__a22o_1 _5420_ (.A1(\mem[11][15] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][15] ),
    .X(_2067_));
 sky130_fd_sc_hd__a2111o_1 _5421_ (.A1(\mem[26][15] ),
    .A2(_1943_),
    .B1(_2065_),
    .C1(_2066_),
    .D1(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__a22o_1 _5422_ (.A1(\mem[16][15] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][15] ),
    .X(_2069_));
 sky130_fd_sc_hd__a221o_1 _5423_ (.A1(\mem[6][15] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][15] ),
    .C1(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__a22o_1 _5424_ (.A1(\mem[28][15] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][15] ),
    .X(_2071_));
 sky130_fd_sc_hd__a221o_1 _5425_ (.A1(\mem[17][15] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][15] ),
    .C1(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__or4_1 _5426_ (.A(_2064_),
    .B(_2068_),
    .C(_2070_),
    .D(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_4 _5427_ (.A(_2073_),
    .X(net56));
 sky130_fd_sc_hd__and3_1 _5428_ (.A(_1822_),
    .B(\mem[24][16] ),
    .C(_1823_),
    .X(_2074_));
 sky130_fd_sc_hd__and3_1 _5429_ (.A(\mem[30][16] ),
    .B(_1854_),
    .C(_2046_),
    .X(_2075_));
 sky130_fd_sc_hd__and3_1 _5430_ (.A(_1856_),
    .B(\mem[27][16] ),
    .C(_1886_),
    .X(_2076_));
 sky130_fd_sc_hd__a2111o_1 _5431_ (.A1(\mem[12][16] ),
    .A2(_1883_),
    .B1(_2074_),
    .C1(_2075_),
    .D1(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__and3_1 _5432_ (.A(_2050_),
    .B(\mem[15][16] ),
    .C(_1889_),
    .X(_2078_));
 sky130_fd_sc_hd__and3b_1 _5433_ (.A_N(_1560_),
    .B(_1599_),
    .C(\mem[13][16] ),
    .X(_2079_));
 sky130_fd_sc_hd__and3_1 _5434_ (.A(_1613_),
    .B(\mem[8][16] ),
    .C(_1861_),
    .X(_2080_));
 sky130_fd_sc_hd__a2111o_1 _5435_ (.A1(\mem[10][16] ),
    .A2(_1926_),
    .B1(_2078_),
    .C1(_2079_),
    .D1(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__inv_2 _5436_ (.A(\mem[3][16] ),
    .Y(_2082_));
 sky130_fd_sc_hd__nor3_1 _5437_ (.A(_2082_),
    .B(_1607_),
    .C(_1688_),
    .Y(_2083_));
 sky130_fd_sc_hd__and4b_1 _5438_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][16] ),
    .D(_1610_),
    .X(_2084_));
 sky130_fd_sc_hd__and3b_1 _5439_ (.A_N(_1556_),
    .B(_2028_),
    .C(\mem[5][16] ),
    .X(_2085_));
 sky130_fd_sc_hd__a2111o_1 _5440_ (.A1(\mem[1][16] ),
    .A2(_1894_),
    .B1(_2083_),
    .C1(_2084_),
    .D1(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_4 _5441_ (.A(_1506_),
    .X(_2087_));
 sky130_fd_sc_hd__and3_1 _5442_ (.A(\mem[18][16] ),
    .B(_1807_),
    .C(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__and3_1 _5443_ (.A(\mem[2][16] ),
    .B(_1838_),
    .C(_1839_),
    .X(_2089_));
 sky130_fd_sc_hd__and3_1 _5444_ (.A(_1903_),
    .B(\mem[23][16] ),
    .C(_1904_),
    .X(_2090_));
 sky130_fd_sc_hd__a2111o_1 _5445_ (.A1(\mem[20][16] ),
    .A2(_1900_),
    .B1(_2088_),
    .C1(_2089_),
    .D1(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__or4_1 _5446_ (.A(_2077_),
    .B(_2081_),
    .C(_2086_),
    .D(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__a22o_1 _5447_ (.A1(\mem[7][16] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][16] ),
    .X(_2093_));
 sky130_fd_sc_hd__a22o_1 _5448_ (.A1(\mem[31][16] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][16] ),
    .X(_2094_));
 sky130_fd_sc_hd__a22o_1 _5449_ (.A1(\mem[11][16] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][16] ),
    .X(_2095_));
 sky130_fd_sc_hd__a2111o_1 _5450_ (.A1(\mem[26][16] ),
    .A2(_1943_),
    .B1(_2093_),
    .C1(_2094_),
    .D1(_2095_),
    .X(_2096_));
 sky130_fd_sc_hd__a22o_1 _5451_ (.A1(\mem[16][16] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][16] ),
    .X(_2097_));
 sky130_fd_sc_hd__a221o_1 _5452_ (.A1(\mem[6][16] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][16] ),
    .C1(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__a22o_1 _5453_ (.A1(\mem[28][16] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][16] ),
    .X(_2099_));
 sky130_fd_sc_hd__a221o_1 _5454_ (.A1(\mem[17][16] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][16] ),
    .C1(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__or4_4 _5455_ (.A(_2092_),
    .B(_2096_),
    .C(_2098_),
    .D(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__clkbuf_1 _5456_ (.A(_2101_),
    .X(net57));
 sky130_fd_sc_hd__and3_1 _5457_ (.A(_1822_),
    .B(\mem[24][17] ),
    .C(_1823_),
    .X(_2102_));
 sky130_fd_sc_hd__and3_1 _5458_ (.A(\mem[30][17] ),
    .B(_1854_),
    .C(_2046_),
    .X(_2103_));
 sky130_fd_sc_hd__and3_1 _5459_ (.A(_1856_),
    .B(\mem[27][17] ),
    .C(_1886_),
    .X(_2104_));
 sky130_fd_sc_hd__a2111o_1 _5460_ (.A1(\mem[12][17] ),
    .A2(_1883_),
    .B1(_2102_),
    .C1(_2103_),
    .D1(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__and3_1 _5461_ (.A(_2050_),
    .B(\mem[15][17] ),
    .C(_1889_),
    .X(_2106_));
 sky130_fd_sc_hd__and3b_1 _5462_ (.A_N(_1560_),
    .B(_1599_),
    .C(\mem[13][17] ),
    .X(_2107_));
 sky130_fd_sc_hd__and3_1 _5463_ (.A(_1613_),
    .B(\mem[8][17] ),
    .C(_1861_),
    .X(_2108_));
 sky130_fd_sc_hd__a2111o_1 _5464_ (.A1(\mem[10][17] ),
    .A2(_1926_),
    .B1(_2106_),
    .C1(_2107_),
    .D1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__inv_2 _5465_ (.A(\mem[3][17] ),
    .Y(_2110_));
 sky130_fd_sc_hd__nor3_1 _5466_ (.A(_2110_),
    .B(_1607_),
    .C(_1688_),
    .Y(_2111_));
 sky130_fd_sc_hd__and4b_1 _5467_ (.A_N(_1536_),
    .B(_1537_),
    .C(\mem[22][17] ),
    .D(_1610_),
    .X(_2112_));
 sky130_fd_sc_hd__and3b_1 _5468_ (.A_N(_1556_),
    .B(_2028_),
    .C(\mem[5][17] ),
    .X(_2113_));
 sky130_fd_sc_hd__a2111o_1 _5469_ (.A1(\mem[1][17] ),
    .A2(_1894_),
    .B1(_2111_),
    .C1(_2112_),
    .D1(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_4 _5470_ (.A(_1503_),
    .X(_2115_));
 sky130_fd_sc_hd__and3_1 _5471_ (.A(\mem[18][17] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2116_));
 sky130_fd_sc_hd__and3_1 _5472_ (.A(\mem[2][17] ),
    .B(_1838_),
    .C(_1839_),
    .X(_2117_));
 sky130_fd_sc_hd__and3_1 _5473_ (.A(_1903_),
    .B(\mem[23][17] ),
    .C(_1904_),
    .X(_2118_));
 sky130_fd_sc_hd__a2111o_1 _5474_ (.A1(\mem[20][17] ),
    .A2(_1900_),
    .B1(_2116_),
    .C1(_2117_),
    .D1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__or4_1 _5475_ (.A(_2105_),
    .B(_2109_),
    .C(_2114_),
    .D(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__a22o_1 _5476_ (.A1(\mem[7][17] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][17] ),
    .X(_2121_));
 sky130_fd_sc_hd__a22o_1 _5477_ (.A1(\mem[31][17] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][17] ),
    .X(_2122_));
 sky130_fd_sc_hd__a22o_1 _5478_ (.A1(\mem[11][17] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][17] ),
    .X(_2123_));
 sky130_fd_sc_hd__a2111o_1 _5479_ (.A1(\mem[26][17] ),
    .A2(_1943_),
    .B1(_2121_),
    .C1(_2122_),
    .D1(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__a22o_1 _5480_ (.A1(\mem[16][17] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][17] ),
    .X(_2125_));
 sky130_fd_sc_hd__a221o_1 _5481_ (.A1(\mem[6][17] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][17] ),
    .C1(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__a22o_1 _5482_ (.A1(\mem[28][17] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][17] ),
    .X(_2127_));
 sky130_fd_sc_hd__a221o_1 _5483_ (.A1(\mem[17][17] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][17] ),
    .C1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__or4_4 _5484_ (.A(_2120_),
    .B(_2124_),
    .C(_2126_),
    .D(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__buf_2 _5485_ (.A(_2129_),
    .X(net58));
 sky130_fd_sc_hd__buf_2 _5486_ (.A(_1519_),
    .X(_2130_));
 sky130_fd_sc_hd__buf_2 _5487_ (.A(_1522_),
    .X(_2131_));
 sky130_fd_sc_hd__and3_1 _5488_ (.A(_2130_),
    .B(\mem[24][18] ),
    .C(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__and3_1 _5489_ (.A(\mem[30][18] ),
    .B(_1854_),
    .C(_2046_),
    .X(_2133_));
 sky130_fd_sc_hd__and3_1 _5490_ (.A(_1856_),
    .B(\mem[27][18] ),
    .C(_1886_),
    .X(_2134_));
 sky130_fd_sc_hd__a2111o_1 _5491_ (.A1(\mem[12][18] ),
    .A2(_1883_),
    .B1(_2132_),
    .C1(_2133_),
    .D1(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__and3_1 _5492_ (.A(_2050_),
    .B(\mem[15][18] ),
    .C(_1889_),
    .X(_2136_));
 sky130_fd_sc_hd__and3b_1 _5493_ (.A_N(_1560_),
    .B(_1599_),
    .C(\mem[13][18] ),
    .X(_2137_));
 sky130_fd_sc_hd__and3_1 _5494_ (.A(_1613_),
    .B(\mem[8][18] ),
    .C(_1861_),
    .X(_2138_));
 sky130_fd_sc_hd__a2111o_1 _5495_ (.A1(\mem[10][18] ),
    .A2(_1926_),
    .B1(_2136_),
    .C1(_2137_),
    .D1(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__and4b_1 _5496_ (.A_N(_1931_),
    .B(_1932_),
    .C(\mem[22][18] ),
    .D(_1507_),
    .X(_2140_));
 sky130_fd_sc_hd__inv_2 _5497_ (.A(\mem[3][18] ),
    .Y(_2141_));
 sky130_fd_sc_hd__nor3_1 _5498_ (.A(_2141_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2142_));
 sky130_fd_sc_hd__and3b_1 _5499_ (.A_N(_1556_),
    .B(_2028_),
    .C(\mem[5][18] ),
    .X(_2143_));
 sky130_fd_sc_hd__a2111o_1 _5500_ (.A1(\mem[1][18] ),
    .A2(_1894_),
    .B1(_2140_),
    .C1(_2142_),
    .D1(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__and3_1 _5501_ (.A(\mem[18][18] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2145_));
 sky130_fd_sc_hd__clkbuf_4 _5502_ (.A(_1504_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_4 _5503_ (.A(_1524_),
    .X(_2147_));
 sky130_fd_sc_hd__and3_1 _5504_ (.A(\mem[2][18] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__and3_1 _5505_ (.A(_1903_),
    .B(\mem[23][18] ),
    .C(_1904_),
    .X(_2149_));
 sky130_fd_sc_hd__a2111o_1 _5506_ (.A1(\mem[20][18] ),
    .A2(_1900_),
    .B1(_2145_),
    .C1(_2148_),
    .D1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__or4_1 _5507_ (.A(_2135_),
    .B(_2139_),
    .C(_2144_),
    .D(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__a22o_1 _5508_ (.A1(\mem[7][18] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][18] ),
    .X(_2152_));
 sky130_fd_sc_hd__a22o_1 _5509_ (.A1(\mem[31][18] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][18] ),
    .X(_2153_));
 sky130_fd_sc_hd__a22o_1 _5510_ (.A1(\mem[11][18] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][18] ),
    .X(_2154_));
 sky130_fd_sc_hd__a2111o_1 _5511_ (.A1(\mem[26][18] ),
    .A2(_1943_),
    .B1(_2152_),
    .C1(_2153_),
    .D1(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__a22o_1 _5512_ (.A1(\mem[16][18] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][18] ),
    .X(_2156_));
 sky130_fd_sc_hd__a221o_1 _5513_ (.A1(\mem[6][18] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][18] ),
    .C1(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__a22o_1 _5514_ (.A1(\mem[28][18] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][18] ),
    .X(_2158_));
 sky130_fd_sc_hd__a221o_1 _5515_ (.A1(\mem[17][18] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][18] ),
    .C1(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__or4_4 _5516_ (.A(_2151_),
    .B(_2155_),
    .C(_2157_),
    .D(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__clkbuf_1 _5517_ (.A(_2160_),
    .X(net59));
 sky130_fd_sc_hd__and3_1 _5518_ (.A(\mem[24][19] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2161_));
 sky130_fd_sc_hd__clkbuf_4 _5519_ (.A(_1509_),
    .X(_2162_));
 sky130_fd_sc_hd__and3_1 _5520_ (.A(\mem[30][19] ),
    .B(_2162_),
    .C(_2046_),
    .X(_2163_));
 sky130_fd_sc_hd__clkbuf_4 _5521_ (.A(_1519_),
    .X(_2164_));
 sky130_fd_sc_hd__and3_1 _5522_ (.A(\mem[27][19] ),
    .B(_2164_),
    .C(_1886_),
    .X(_2165_));
 sky130_fd_sc_hd__a2111o_1 _5523_ (.A1(\mem[12][19] ),
    .A2(_1883_),
    .B1(_2161_),
    .C1(_2163_),
    .D1(_2165_),
    .X(_2166_));
 sky130_fd_sc_hd__and3_1 _5524_ (.A(\mem[15][19] ),
    .B(_2050_),
    .C(_1889_),
    .X(_2167_));
 sky130_fd_sc_hd__clkbuf_4 _5525_ (.A(_1499_),
    .X(_2168_));
 sky130_fd_sc_hd__nor3b_1 _5526_ (.A(_2168_),
    .B(_1561_),
    .C_N(\mem[13][19] ),
    .Y(_2169_));
 sky130_fd_sc_hd__clkbuf_4 _5527_ (.A(_1522_),
    .X(_2170_));
 sky130_fd_sc_hd__and3_1 _5528_ (.A(\mem[8][19] ),
    .B(_2028_),
    .C(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__a2111o_1 _5529_ (.A1(\mem[10][19] ),
    .A2(_1926_),
    .B1(_2167_),
    .C1(_2169_),
    .D1(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__nor3_1 _5530_ (.A(_1031_),
    .B(_1607_),
    .C(_1688_),
    .Y(_2173_));
 sky130_fd_sc_hd__clkbuf_4 _5531_ (.A(_1506_),
    .X(_2174_));
 sky130_fd_sc_hd__and4b_1 _5532_ (.A_N(_1536_),
    .B(_1537_),
    .C(_2174_),
    .D(\mem[22][19] ),
    .X(_2175_));
 sky130_fd_sc_hd__nor3b_1 _5533_ (.A(_1514_),
    .B(_1557_),
    .C_N(\mem[5][19] ),
    .Y(_2176_));
 sky130_fd_sc_hd__a2111o_1 _5534_ (.A1(\mem[1][19] ),
    .A2(_1894_),
    .B1(_2173_),
    .C1(_2175_),
    .D1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__and3_1 _5535_ (.A(\mem[18][19] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2178_));
 sky130_fd_sc_hd__and3_1 _5536_ (.A(\mem[2][19] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2179_));
 sky130_fd_sc_hd__and3_1 _5537_ (.A(\mem[23][19] ),
    .B(_1903_),
    .C(_1904_),
    .X(_2180_));
 sky130_fd_sc_hd__a2111o_1 _5538_ (.A1(\mem[20][19] ),
    .A2(_1900_),
    .B1(_2178_),
    .C1(_2179_),
    .D1(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__or4_1 _5539_ (.A(_2166_),
    .B(_2172_),
    .C(_2177_),
    .D(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__a22o_1 _5540_ (.A1(\mem[7][19] ),
    .A2(_1908_),
    .B1(_1909_),
    .B2(\mem[9][19] ),
    .X(_2183_));
 sky130_fd_sc_hd__a22o_1 _5541_ (.A1(\mem[31][19] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][19] ),
    .X(_2184_));
 sky130_fd_sc_hd__a22o_1 _5542_ (.A1(\mem[11][19] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][19] ),
    .X(_2185_));
 sky130_fd_sc_hd__a2111o_1 _5543_ (.A1(\mem[26][19] ),
    .A2(_1943_),
    .B1(_2183_),
    .C1(_2184_),
    .D1(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__a22o_1 _5544_ (.A1(\mem[16][19] ),
    .A2(_1914_),
    .B1(_1915_),
    .B2(\mem[19][19] ),
    .X(_2187_));
 sky130_fd_sc_hd__a221o_1 _5545_ (.A1(\mem[6][19] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][19] ),
    .C1(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__a22o_1 _5546_ (.A1(\mem[28][19] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][19] ),
    .X(_2189_));
 sky130_fd_sc_hd__a221o_1 _5547_ (.A1(\mem[17][19] ),
    .A2(_1918_),
    .B1(_1956_),
    .B2(\mem[21][19] ),
    .C1(_2189_),
    .X(_2190_));
 sky130_fd_sc_hd__or4_1 _5548_ (.A(_2182_),
    .B(_2186_),
    .C(_2188_),
    .D(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__buf_6 _5549_ (.A(_2191_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 _5550_ (.A(_1511_),
    .X(_2192_));
 sky130_fd_sc_hd__and3_1 _5551_ (.A(\mem[24][20] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2193_));
 sky130_fd_sc_hd__and3_1 _5552_ (.A(\mem[30][20] ),
    .B(_2162_),
    .C(_2046_),
    .X(_2194_));
 sky130_fd_sc_hd__buf_2 _5553_ (.A(_1497_),
    .X(_2195_));
 sky130_fd_sc_hd__and3_1 _5554_ (.A(\mem[27][20] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__a2111o_1 _5555_ (.A1(\mem[12][20] ),
    .A2(_2192_),
    .B1(_2193_),
    .C1(_2194_),
    .D1(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__buf_2 _5556_ (.A(_1500_),
    .X(_2198_));
 sky130_fd_sc_hd__and3_1 _5557_ (.A(\mem[15][20] ),
    .B(_2050_),
    .C(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__nor3b_1 _5558_ (.A(_2168_),
    .B(_1561_),
    .C_N(\mem[13][20] ),
    .Y(_2200_));
 sky130_fd_sc_hd__and3_1 _5559_ (.A(\mem[8][20] ),
    .B(_2028_),
    .C(_2170_),
    .X(_2201_));
 sky130_fd_sc_hd__a2111o_1 _5560_ (.A1(\mem[10][20] ),
    .A2(_1926_),
    .B1(_2199_),
    .C1(_2200_),
    .D1(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_4 _5561_ (.A(_1550_),
    .X(_2203_));
 sky130_fd_sc_hd__nor3_1 _5562_ (.A(_1113_),
    .B(_1607_),
    .C(_1688_),
    .Y(_2204_));
 sky130_fd_sc_hd__and4b_1 _5563_ (.A_N(_1536_),
    .B(_1537_),
    .C(_2174_),
    .D(\mem[22][20] ),
    .X(_2205_));
 sky130_fd_sc_hd__nor3b_1 _5564_ (.A(_1514_),
    .B(_1557_),
    .C_N(\mem[5][20] ),
    .Y(_2206_));
 sky130_fd_sc_hd__a2111o_1 _5565_ (.A1(\mem[1][20] ),
    .A2(_2203_),
    .B1(_2204_),
    .C1(_2205_),
    .D1(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_4 _5566_ (.A(_1541_),
    .X(_2208_));
 sky130_fd_sc_hd__and3_1 _5567_ (.A(\mem[18][20] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2209_));
 sky130_fd_sc_hd__and3_1 _5568_ (.A(\mem[2][20] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2210_));
 sky130_fd_sc_hd__buf_2 _5569_ (.A(_1519_),
    .X(_2211_));
 sky130_fd_sc_hd__buf_2 _5570_ (.A(_1564_),
    .X(_2212_));
 sky130_fd_sc_hd__and3_1 _5571_ (.A(\mem[23][20] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__a2111o_1 _5572_ (.A1(\mem[20][20] ),
    .A2(_2208_),
    .B1(_2209_),
    .C1(_2210_),
    .D1(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__or4_1 _5573_ (.A(_2197_),
    .B(_2202_),
    .C(_2207_),
    .D(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__clkbuf_4 _5574_ (.A(_1565_),
    .X(_2216_));
 sky130_fd_sc_hd__clkbuf_4 _5575_ (.A(_1571_),
    .X(_2217_));
 sky130_fd_sc_hd__a22o_1 _5576_ (.A1(\mem[7][20] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][20] ),
    .X(_2218_));
 sky130_fd_sc_hd__a22o_1 _5577_ (.A1(\mem[31][20] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(\mem[25][20] ),
    .X(_2219_));
 sky130_fd_sc_hd__a22o_1 _5578_ (.A1(\mem[11][20] ),
    .A2(_1948_),
    .B1(_1949_),
    .B2(\mem[14][20] ),
    .X(_2220_));
 sky130_fd_sc_hd__a2111o_1 _5579_ (.A1(\mem[26][20] ),
    .A2(_1943_),
    .B1(_2218_),
    .C1(_2219_),
    .D1(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__clkbuf_4 _5580_ (.A(_1546_),
    .X(_2222_));
 sky130_fd_sc_hd__clkbuf_4 _5581_ (.A(_1580_),
    .X(_2223_));
 sky130_fd_sc_hd__a22o_1 _5582_ (.A1(\mem[16][20] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][20] ),
    .X(_2224_));
 sky130_fd_sc_hd__a221o_1 _5583_ (.A1(\mem[6][20] ),
    .A2(_1952_),
    .B1(_1953_),
    .B2(\mem[4][20] ),
    .C1(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__buf_4 _5584_ (.A(_1530_),
    .X(_2226_));
 sky130_fd_sc_hd__a22o_1 _5585_ (.A1(\mem[28][20] ),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\mem[29][20] ),
    .X(_2227_));
 sky130_fd_sc_hd__a221o_1 _5586_ (.A1(\mem[17][20] ),
    .A2(_2226_),
    .B1(_1956_),
    .B2(\mem[21][20] ),
    .C1(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__or4_4 _5587_ (.A(_2215_),
    .B(_2221_),
    .C(_2225_),
    .D(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_1 _5588_ (.A(_2229_),
    .X(net62));
 sky130_fd_sc_hd__and3_1 _5589_ (.A(\mem[24][21] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2230_));
 sky130_fd_sc_hd__and3_1 _5590_ (.A(\mem[30][21] ),
    .B(_2162_),
    .C(_2046_),
    .X(_2231_));
 sky130_fd_sc_hd__and3_1 _5591_ (.A(\mem[27][21] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2232_));
 sky130_fd_sc_hd__a2111o_1 _5592_ (.A1(\mem[12][21] ),
    .A2(_2192_),
    .B1(_2230_),
    .C1(_2231_),
    .D1(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__clkbuf_4 _5593_ (.A(_1597_),
    .X(_2234_));
 sky130_fd_sc_hd__and3_1 _5594_ (.A(\mem[15][21] ),
    .B(_2050_),
    .C(_2198_),
    .X(_2235_));
 sky130_fd_sc_hd__clkbuf_4 _5595_ (.A(_1499_),
    .X(_2236_));
 sky130_fd_sc_hd__nor3b_1 _5596_ (.A(_2236_),
    .B(_1561_),
    .C_N(\mem[13][21] ),
    .Y(_2237_));
 sky130_fd_sc_hd__and3_1 _5597_ (.A(\mem[8][21] ),
    .B(_2028_),
    .C(_2170_),
    .X(_2238_));
 sky130_fd_sc_hd__a2111o_1 _5598_ (.A1(\mem[10][21] ),
    .A2(_2234_),
    .B1(_2235_),
    .C1(_2237_),
    .D1(_2238_),
    .X(_2239_));
 sky130_fd_sc_hd__and4b_1 _5599_ (.A_N(_1931_),
    .B(_1932_),
    .C(_1610_),
    .D(\mem[22][21] ),
    .X(_2240_));
 sky130_fd_sc_hd__nor3_1 _5600_ (.A(_1150_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2241_));
 sky130_fd_sc_hd__nor3b_1 _5601_ (.A(_1514_),
    .B(_1557_),
    .C_N(\mem[5][21] ),
    .Y(_2242_));
 sky130_fd_sc_hd__a2111o_1 _5602_ (.A1(\mem[1][21] ),
    .A2(_2203_),
    .B1(_2240_),
    .C1(_2241_),
    .D1(_2242_),
    .X(_2243_));
 sky130_fd_sc_hd__and3_1 _5603_ (.A(\mem[18][21] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2244_));
 sky130_fd_sc_hd__and3_1 _5604_ (.A(\mem[2][21] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2245_));
 sky130_fd_sc_hd__and3_1 _5605_ (.A(\mem[23][21] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2246_));
 sky130_fd_sc_hd__a2111o_1 _5606_ (.A1(\mem[20][21] ),
    .A2(_2208_),
    .B1(_2244_),
    .C1(_2245_),
    .D1(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__or4_1 _5607_ (.A(_2233_),
    .B(_2239_),
    .C(_2243_),
    .D(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__clkbuf_4 _5608_ (.A(_1623_),
    .X(_2249_));
 sky130_fd_sc_hd__a22o_1 _5609_ (.A1(\mem[7][21] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][21] ),
    .X(_2250_));
 sky130_fd_sc_hd__clkbuf_4 _5610_ (.A(_1501_),
    .X(_2251_));
 sky130_fd_sc_hd__clkbuf_4 _5611_ (.A(_1520_),
    .X(_2252_));
 sky130_fd_sc_hd__a22o_1 _5612_ (.A1(\mem[31][21] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][21] ),
    .X(_2253_));
 sky130_fd_sc_hd__clkbuf_4 _5613_ (.A(_1498_),
    .X(_2254_));
 sky130_fd_sc_hd__clkbuf_4 _5614_ (.A(_1525_),
    .X(_2255_));
 sky130_fd_sc_hd__a22o_1 _5615_ (.A1(\mem[11][21] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][21] ),
    .X(_2256_));
 sky130_fd_sc_hd__a2111o_1 _5616_ (.A1(\mem[26][21] ),
    .A2(_2249_),
    .B1(_2250_),
    .C1(_2253_),
    .D1(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__clkbuf_4 _5617_ (.A(_1539_),
    .X(_2258_));
 sky130_fd_sc_hd__clkbuf_4 _5618_ (.A(_1554_),
    .X(_2259_));
 sky130_fd_sc_hd__a22o_1 _5619_ (.A1(\mem[16][21] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][21] ),
    .X(_2260_));
 sky130_fd_sc_hd__a221o_1 _5620_ (.A1(\mem[6][21] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][21] ),
    .C1(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__buf_4 _5621_ (.A(_1637_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_4 _5622_ (.A(_1639_),
    .X(_2263_));
 sky130_fd_sc_hd__clkbuf_4 _5623_ (.A(_1641_),
    .X(_2264_));
 sky130_fd_sc_hd__a22o_1 _5624_ (.A1(\mem[28][21] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][21] ),
    .X(_2265_));
 sky130_fd_sc_hd__a221o_1 _5625_ (.A1(\mem[17][21] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][21] ),
    .C1(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__or4_4 _5626_ (.A(_2248_),
    .B(_2257_),
    .C(_2261_),
    .D(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__buf_4 _5627_ (.A(_2267_),
    .X(net63));
 sky130_fd_sc_hd__and3_1 _5628_ (.A(\mem[24][22] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2268_));
 sky130_fd_sc_hd__and3_1 _5629_ (.A(\mem[30][22] ),
    .B(_2162_),
    .C(_2046_),
    .X(_2269_));
 sky130_fd_sc_hd__and3_1 _5630_ (.A(\mem[27][22] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2270_));
 sky130_fd_sc_hd__a2111o_1 _5631_ (.A1(\mem[12][22] ),
    .A2(_2192_),
    .B1(_2268_),
    .C1(_2269_),
    .D1(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__and3_1 _5632_ (.A(\mem[15][22] ),
    .B(_2050_),
    .C(_2198_),
    .X(_2272_));
 sky130_fd_sc_hd__nor3b_1 _5633_ (.A(_2236_),
    .B(_1561_),
    .C_N(\mem[13][22] ),
    .Y(_2273_));
 sky130_fd_sc_hd__and3_1 _5634_ (.A(\mem[8][22] ),
    .B(_2028_),
    .C(_2170_),
    .X(_2274_));
 sky130_fd_sc_hd__a2111o_1 _5635_ (.A1(\mem[10][22] ),
    .A2(_2234_),
    .B1(_2272_),
    .C1(_2273_),
    .D1(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__and4b_1 _5636_ (.A_N(_1931_),
    .B(_1932_),
    .C(_1657_),
    .D(\mem[22][22] ),
    .X(_2276_));
 sky130_fd_sc_hd__nor3_1 _5637_ (.A(_1179_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2277_));
 sky130_fd_sc_hd__nor3b_1 _5638_ (.A(_1514_),
    .B(_1557_),
    .C_N(\mem[5][22] ),
    .Y(_2278_));
 sky130_fd_sc_hd__a2111o_1 _5639_ (.A1(\mem[1][22] ),
    .A2(_2203_),
    .B1(_2276_),
    .C1(_2277_),
    .D1(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__and3_1 _5640_ (.A(\mem[18][22] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2280_));
 sky130_fd_sc_hd__and3_1 _5641_ (.A(\mem[2][22] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2281_));
 sky130_fd_sc_hd__and3_1 _5642_ (.A(\mem[23][22] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2282_));
 sky130_fd_sc_hd__a2111o_1 _5643_ (.A1(\mem[20][22] ),
    .A2(_2208_),
    .B1(_2280_),
    .C1(_2281_),
    .D1(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__or4_1 _5644_ (.A(_2271_),
    .B(_2275_),
    .C(_2279_),
    .D(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__a22o_1 _5645_ (.A1(\mem[7][22] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][22] ),
    .X(_2285_));
 sky130_fd_sc_hd__a22o_1 _5646_ (.A1(\mem[31][22] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][22] ),
    .X(_2286_));
 sky130_fd_sc_hd__a22o_1 _5647_ (.A1(\mem[11][22] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][22] ),
    .X(_2287_));
 sky130_fd_sc_hd__a2111o_1 _5648_ (.A1(\mem[26][22] ),
    .A2(_2249_),
    .B1(_2285_),
    .C1(_2286_),
    .D1(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__a22o_1 _5649_ (.A1(\mem[16][22] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][22] ),
    .X(_2289_));
 sky130_fd_sc_hd__a221o_1 _5650_ (.A1(\mem[6][22] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][22] ),
    .C1(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__a22o_1 _5651_ (.A1(\mem[28][22] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][22] ),
    .X(_2291_));
 sky130_fd_sc_hd__a221o_1 _5652_ (.A1(\mem[17][22] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][22] ),
    .C1(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__or4_4 _5653_ (.A(_2284_),
    .B(_2288_),
    .C(_2290_),
    .D(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__clkbuf_1 _5654_ (.A(_2293_),
    .X(net64));
 sky130_fd_sc_hd__and3_1 _5655_ (.A(\mem[24][23] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2294_));
 sky130_fd_sc_hd__and3_1 _5656_ (.A(\mem[30][23] ),
    .B(_2162_),
    .C(_2046_),
    .X(_2295_));
 sky130_fd_sc_hd__and3_1 _5657_ (.A(\mem[27][23] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2296_));
 sky130_fd_sc_hd__a2111o_1 _5658_ (.A1(\mem[12][23] ),
    .A2(_2192_),
    .B1(_2294_),
    .C1(_2295_),
    .D1(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__and3_1 _5659_ (.A(\mem[15][23] ),
    .B(_2050_),
    .C(_2198_),
    .X(_2298_));
 sky130_fd_sc_hd__nor3b_1 _5660_ (.A(_2236_),
    .B(_1561_),
    .C_N(\mem[13][23] ),
    .Y(_2299_));
 sky130_fd_sc_hd__and3_1 _5661_ (.A(\mem[8][23] ),
    .B(_2028_),
    .C(_2170_),
    .X(_2300_));
 sky130_fd_sc_hd__a2111o_1 _5662_ (.A1(\mem[10][23] ),
    .A2(_2234_),
    .B1(_2298_),
    .C1(_2299_),
    .D1(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__and4b_1 _5663_ (.A_N(_1931_),
    .B(_1932_),
    .C(_1657_),
    .D(\mem[22][23] ),
    .X(_2302_));
 sky130_fd_sc_hd__nor3_1 _5664_ (.A(_1210_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2303_));
 sky130_fd_sc_hd__nor3b_1 _5665_ (.A(_1514_),
    .B(_1557_),
    .C_N(\mem[5][23] ),
    .Y(_2304_));
 sky130_fd_sc_hd__a2111o_1 _5666_ (.A1(\mem[1][23] ),
    .A2(_2203_),
    .B1(_2302_),
    .C1(_2303_),
    .D1(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__and3_1 _5667_ (.A(\mem[18][23] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2306_));
 sky130_fd_sc_hd__and3_1 _5668_ (.A(\mem[2][23] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2307_));
 sky130_fd_sc_hd__and3_1 _5669_ (.A(\mem[23][23] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2308_));
 sky130_fd_sc_hd__a2111o_1 _5670_ (.A1(\mem[20][23] ),
    .A2(_2208_),
    .B1(_2306_),
    .C1(_2307_),
    .D1(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__or4_1 _5671_ (.A(_2297_),
    .B(_2301_),
    .C(_2305_),
    .D(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__a22o_1 _5672_ (.A1(\mem[7][23] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][23] ),
    .X(_2311_));
 sky130_fd_sc_hd__a22o_1 _5673_ (.A1(\mem[31][23] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][23] ),
    .X(_2312_));
 sky130_fd_sc_hd__a22o_1 _5674_ (.A1(\mem[11][23] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][23] ),
    .X(_2313_));
 sky130_fd_sc_hd__a2111o_1 _5675_ (.A1(\mem[26][23] ),
    .A2(_2249_),
    .B1(_2311_),
    .C1(_2312_),
    .D1(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__a22o_1 _5676_ (.A1(\mem[16][23] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][23] ),
    .X(_2315_));
 sky130_fd_sc_hd__a221o_1 _5677_ (.A1(\mem[6][23] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][23] ),
    .C1(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__a22o_1 _5678_ (.A1(\mem[28][23] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][23] ),
    .X(_2317_));
 sky130_fd_sc_hd__a221o_1 _5679_ (.A1(\mem[17][23] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][23] ),
    .C1(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__or4_1 _5680_ (.A(_2310_),
    .B(_2314_),
    .C(_2316_),
    .D(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__buf_4 _5681_ (.A(_2319_),
    .X(net65));
 sky130_fd_sc_hd__and3_1 _5682_ (.A(\mem[24][24] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2320_));
 sky130_fd_sc_hd__and3_1 _5683_ (.A(\mem[30][24] ),
    .B(_2162_),
    .C(_2046_),
    .X(_2321_));
 sky130_fd_sc_hd__and3_1 _5684_ (.A(\mem[27][24] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2322_));
 sky130_fd_sc_hd__a2111o_1 _5685_ (.A1(\mem[12][24] ),
    .A2(_2192_),
    .B1(_2320_),
    .C1(_2321_),
    .D1(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__and3_1 _5686_ (.A(\mem[15][24] ),
    .B(_2050_),
    .C(_2198_),
    .X(_2324_));
 sky130_fd_sc_hd__nor3b_1 _5687_ (.A(_2236_),
    .B(_1561_),
    .C_N(\mem[13][24] ),
    .Y(_2325_));
 sky130_fd_sc_hd__and3_1 _5688_ (.A(\mem[8][24] ),
    .B(_1602_),
    .C(_2170_),
    .X(_2326_));
 sky130_fd_sc_hd__a2111o_1 _5689_ (.A1(\mem[10][24] ),
    .A2(_2234_),
    .B1(_2324_),
    .C1(_2325_),
    .D1(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__and4b_1 _5690_ (.A_N(_1931_),
    .B(_1932_),
    .C(_1657_),
    .D(\mem[22][24] ),
    .X(_2328_));
 sky130_fd_sc_hd__nor3_1 _5691_ (.A(_1240_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2329_));
 sky130_fd_sc_hd__nor3b_1 _5692_ (.A(_2168_),
    .B(_1557_),
    .C_N(\mem[5][24] ),
    .Y(_2330_));
 sky130_fd_sc_hd__a2111o_1 _5693_ (.A1(\mem[1][24] ),
    .A2(_2203_),
    .B1(_2328_),
    .C1(_2329_),
    .D1(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__and3_1 _5694_ (.A(\mem[18][24] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2332_));
 sky130_fd_sc_hd__and3_1 _5695_ (.A(\mem[2][24] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2333_));
 sky130_fd_sc_hd__and3_1 _5696_ (.A(\mem[23][24] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2334_));
 sky130_fd_sc_hd__a2111o_1 _5697_ (.A1(\mem[20][24] ),
    .A2(_2208_),
    .B1(_2332_),
    .C1(_2333_),
    .D1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__or4_1 _5698_ (.A(_2323_),
    .B(_2327_),
    .C(_2331_),
    .D(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__a22o_1 _5699_ (.A1(\mem[7][24] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][24] ),
    .X(_2337_));
 sky130_fd_sc_hd__a22o_1 _5700_ (.A1(\mem[31][24] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][24] ),
    .X(_2338_));
 sky130_fd_sc_hd__a22o_1 _5701_ (.A1(\mem[11][24] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][24] ),
    .X(_2339_));
 sky130_fd_sc_hd__a2111o_1 _5702_ (.A1(\mem[26][24] ),
    .A2(_2249_),
    .B1(_2337_),
    .C1(_2338_),
    .D1(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__a22o_1 _5703_ (.A1(\mem[16][24] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][24] ),
    .X(_2341_));
 sky130_fd_sc_hd__a221o_1 _5704_ (.A1(\mem[6][24] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][24] ),
    .C1(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__a22o_1 _5705_ (.A1(\mem[28][24] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][24] ),
    .X(_2343_));
 sky130_fd_sc_hd__a221o_1 _5706_ (.A1(\mem[17][24] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][24] ),
    .C1(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__or4_4 _5707_ (.A(_2336_),
    .B(_2340_),
    .C(_2342_),
    .D(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__buf_4 _5708_ (.A(_2345_),
    .X(net66));
 sky130_fd_sc_hd__and3_1 _5709_ (.A(\mem[24][25] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2346_));
 sky130_fd_sc_hd__and3_1 _5710_ (.A(\mem[30][25] ),
    .B(_2162_),
    .C(_2174_),
    .X(_2347_));
 sky130_fd_sc_hd__and3_1 _5711_ (.A(\mem[27][25] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2348_));
 sky130_fd_sc_hd__a2111o_1 _5712_ (.A1(\mem[12][25] ),
    .A2(_2192_),
    .B1(_2346_),
    .C1(_2347_),
    .D1(_2348_),
    .X(_2349_));
 sky130_fd_sc_hd__and3_1 _5713_ (.A(\mem[15][25] ),
    .B(_1494_),
    .C(_2198_),
    .X(_2350_));
 sky130_fd_sc_hd__nor3b_1 _5714_ (.A(_2236_),
    .B(_1561_),
    .C_N(\mem[13][25] ),
    .Y(_2351_));
 sky130_fd_sc_hd__and3_1 _5715_ (.A(\mem[8][25] ),
    .B(_1602_),
    .C(_2170_),
    .X(_2352_));
 sky130_fd_sc_hd__a2111o_1 _5716_ (.A1(\mem[10][25] ),
    .A2(_2234_),
    .B1(_2350_),
    .C1(_2351_),
    .D1(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__nor3_1 _5717_ (.A(_1269_),
    .B(_1607_),
    .C(_1688_),
    .Y(_2354_));
 sky130_fd_sc_hd__and4b_1 _5718_ (.A_N(_1655_),
    .B(_1656_),
    .C(_2174_),
    .D(\mem[22][25] ),
    .X(_2355_));
 sky130_fd_sc_hd__nor3b_1 _5719_ (.A(_2168_),
    .B(_1557_),
    .C_N(\mem[5][25] ),
    .Y(_2356_));
 sky130_fd_sc_hd__a2111o_1 _5720_ (.A1(\mem[1][25] ),
    .A2(_2203_),
    .B1(_2354_),
    .C1(_2355_),
    .D1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__and3_1 _5721_ (.A(\mem[18][25] ),
    .B(_2115_),
    .C(_2087_),
    .X(_2358_));
 sky130_fd_sc_hd__and3_1 _5722_ (.A(\mem[2][25] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2359_));
 sky130_fd_sc_hd__and3_1 _5723_ (.A(\mem[23][25] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2360_));
 sky130_fd_sc_hd__a2111o_1 _5724_ (.A1(\mem[20][25] ),
    .A2(_2208_),
    .B1(_2358_),
    .C1(_2359_),
    .D1(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__or4_1 _5725_ (.A(_2349_),
    .B(_2353_),
    .C(_2357_),
    .D(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__a22o_1 _5726_ (.A1(\mem[7][25] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][25] ),
    .X(_2363_));
 sky130_fd_sc_hd__a22o_1 _5727_ (.A1(\mem[31][25] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][25] ),
    .X(_2364_));
 sky130_fd_sc_hd__a22o_1 _5728_ (.A1(\mem[11][25] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][25] ),
    .X(_2365_));
 sky130_fd_sc_hd__a2111o_1 _5729_ (.A1(\mem[26][25] ),
    .A2(_2249_),
    .B1(_2363_),
    .C1(_2364_),
    .D1(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__a22o_1 _5730_ (.A1(\mem[16][25] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][25] ),
    .X(_2367_));
 sky130_fd_sc_hd__a221o_1 _5731_ (.A1(\mem[6][25] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][25] ),
    .C1(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__a22o_1 _5732_ (.A1(\mem[28][25] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][25] ),
    .X(_2369_));
 sky130_fd_sc_hd__a221o_1 _5733_ (.A1(\mem[17][25] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][25] ),
    .C1(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__or4_2 _5734_ (.A(_2362_),
    .B(_2366_),
    .C(_2368_),
    .D(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__clkbuf_4 _5735_ (.A(_2371_),
    .X(net67));
 sky130_fd_sc_hd__and3_1 _5736_ (.A(\mem[24][26] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2372_));
 sky130_fd_sc_hd__and3_1 _5737_ (.A(\mem[30][26] ),
    .B(_2162_),
    .C(_2174_),
    .X(_2373_));
 sky130_fd_sc_hd__and3_1 _5738_ (.A(\mem[27][26] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2374_));
 sky130_fd_sc_hd__a2111o_1 _5739_ (.A1(\mem[12][26] ),
    .A2(_2192_),
    .B1(_2372_),
    .C1(_2373_),
    .D1(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__and3_1 _5740_ (.A(\mem[15][26] ),
    .B(_1494_),
    .C(_2198_),
    .X(_2376_));
 sky130_fd_sc_hd__nor3b_1 _5741_ (.A(_2236_),
    .B(_1561_),
    .C_N(\mem[13][26] ),
    .Y(_2377_));
 sky130_fd_sc_hd__and3_1 _5742_ (.A(\mem[8][26] ),
    .B(_1602_),
    .C(_2170_),
    .X(_2378_));
 sky130_fd_sc_hd__a2111o_1 _5743_ (.A1(\mem[10][26] ),
    .A2(_2234_),
    .B1(_2376_),
    .C1(_2377_),
    .D1(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__and4b_1 _5744_ (.A_N(_1517_),
    .B(_1516_),
    .C(_1657_),
    .D(\mem[22][26] ),
    .X(_2380_));
 sky130_fd_sc_hd__nor3_1 _5745_ (.A(_1299_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2381_));
 sky130_fd_sc_hd__nor3b_1 _5746_ (.A(_2168_),
    .B(_1612_),
    .C_N(\mem[5][26] ),
    .Y(_2382_));
 sky130_fd_sc_hd__a2111o_1 _5747_ (.A1(\mem[1][26] ),
    .A2(_2203_),
    .B1(_2380_),
    .C1(_2381_),
    .D1(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__and3_1 _5748_ (.A(\mem[18][26] ),
    .B(_2115_),
    .C(_1592_),
    .X(_2384_));
 sky130_fd_sc_hd__and3_1 _5749_ (.A(\mem[2][26] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2385_));
 sky130_fd_sc_hd__and3_1 _5750_ (.A(\mem[23][26] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2386_));
 sky130_fd_sc_hd__a2111o_1 _5751_ (.A1(\mem[20][26] ),
    .A2(_2208_),
    .B1(_2384_),
    .C1(_2385_),
    .D1(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__or4_1 _5752_ (.A(_2375_),
    .B(_2379_),
    .C(_2383_),
    .D(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__a22o_1 _5753_ (.A1(\mem[7][26] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][26] ),
    .X(_2389_));
 sky130_fd_sc_hd__a22o_1 _5754_ (.A1(\mem[31][26] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][26] ),
    .X(_2390_));
 sky130_fd_sc_hd__a22o_1 _5755_ (.A1(\mem[11][26] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][26] ),
    .X(_2391_));
 sky130_fd_sc_hd__a2111o_1 _5756_ (.A1(\mem[26][26] ),
    .A2(_2249_),
    .B1(_2389_),
    .C1(_2390_),
    .D1(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__a22o_1 _5757_ (.A1(\mem[16][26] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][26] ),
    .X(_2393_));
 sky130_fd_sc_hd__a221o_1 _5758_ (.A1(\mem[6][26] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][26] ),
    .C1(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__a22o_1 _5759_ (.A1(\mem[28][26] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][26] ),
    .X(_2395_));
 sky130_fd_sc_hd__a221o_1 _5760_ (.A1(\mem[17][26] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][26] ),
    .C1(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__or4_2 _5761_ (.A(_2388_),
    .B(_2392_),
    .C(_2394_),
    .D(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__buf_4 _5762_ (.A(_2397_),
    .X(net68));
 sky130_fd_sc_hd__and3_1 _5763_ (.A(\mem[24][27] ),
    .B(_2130_),
    .C(_2131_),
    .X(_2398_));
 sky130_fd_sc_hd__and3_1 _5764_ (.A(\mem[30][27] ),
    .B(_2162_),
    .C(_2174_),
    .X(_2399_));
 sky130_fd_sc_hd__and3_1 _5765_ (.A(\mem[27][27] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2400_));
 sky130_fd_sc_hd__a2111o_1 _5766_ (.A1(\mem[12][27] ),
    .A2(_2192_),
    .B1(_2398_),
    .C1(_2399_),
    .D1(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__and3_1 _5767_ (.A(\mem[15][27] ),
    .B(_1494_),
    .C(_2198_),
    .X(_2402_));
 sky130_fd_sc_hd__nor3b_1 _5768_ (.A(_2236_),
    .B(_1601_),
    .C_N(\mem[13][27] ),
    .Y(_2403_));
 sky130_fd_sc_hd__and3_1 _5769_ (.A(\mem[8][27] ),
    .B(_1602_),
    .C(_2170_),
    .X(_2404_));
 sky130_fd_sc_hd__a2111o_1 _5770_ (.A1(\mem[10][27] ),
    .A2(_2234_),
    .B1(_2402_),
    .C1(_2403_),
    .D1(_2404_),
    .X(_2405_));
 sky130_fd_sc_hd__and4b_1 _5771_ (.A_N(_1517_),
    .B(_1516_),
    .C(_1657_),
    .D(\mem[22][27] ),
    .X(_2406_));
 sky130_fd_sc_hd__nor3_1 _5772_ (.A(_1330_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2407_));
 sky130_fd_sc_hd__nor3b_1 _5773_ (.A(_2168_),
    .B(_1612_),
    .C_N(\mem[5][27] ),
    .Y(_2408_));
 sky130_fd_sc_hd__a2111o_1 _5774_ (.A1(\mem[1][27] ),
    .A2(_2203_),
    .B1(_2406_),
    .C1(_2407_),
    .D1(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__and3_1 _5775_ (.A(\mem[18][27] ),
    .B(_1504_),
    .C(_1592_),
    .X(_2410_));
 sky130_fd_sc_hd__and3_1 _5776_ (.A(\mem[2][27] ),
    .B(_2146_),
    .C(_2147_),
    .X(_2411_));
 sky130_fd_sc_hd__and3_1 _5777_ (.A(\mem[23][27] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2412_));
 sky130_fd_sc_hd__a2111o_1 _5778_ (.A1(\mem[20][27] ),
    .A2(_2208_),
    .B1(_2410_),
    .C1(_2411_),
    .D1(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__or4_1 _5779_ (.A(_2401_),
    .B(_2405_),
    .C(_2409_),
    .D(_2413_),
    .X(_2414_));
 sky130_fd_sc_hd__a22o_1 _5780_ (.A1(\mem[7][27] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][27] ),
    .X(_2415_));
 sky130_fd_sc_hd__a22o_1 _5781_ (.A1(\mem[31][27] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][27] ),
    .X(_2416_));
 sky130_fd_sc_hd__a22o_1 _5782_ (.A1(\mem[11][27] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][27] ),
    .X(_2417_));
 sky130_fd_sc_hd__a2111o_1 _5783_ (.A1(\mem[26][27] ),
    .A2(_2249_),
    .B1(_2415_),
    .C1(_2416_),
    .D1(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__a22o_1 _5784_ (.A1(\mem[16][27] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][27] ),
    .X(_2419_));
 sky130_fd_sc_hd__a221o_1 _5785_ (.A1(\mem[6][27] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][27] ),
    .C1(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__a22o_1 _5786_ (.A1(\mem[28][27] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][27] ),
    .X(_2421_));
 sky130_fd_sc_hd__a221o_1 _5787_ (.A1(\mem[17][27] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][27] ),
    .C1(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__or4_4 _5788_ (.A(_2414_),
    .B(_2418_),
    .C(_2420_),
    .D(_2422_),
    .X(_2423_));
 sky130_fd_sc_hd__clkbuf_1 _5789_ (.A(_2423_),
    .X(net69));
 sky130_fd_sc_hd__and3_1 _5790_ (.A(\mem[24][28] ),
    .B(_1499_),
    .C(_1522_),
    .X(_2424_));
 sky130_fd_sc_hd__and3_1 _5791_ (.A(\mem[30][28] ),
    .B(_2162_),
    .C(_2174_),
    .X(_2425_));
 sky130_fd_sc_hd__and3_1 _5792_ (.A(\mem[27][28] ),
    .B(_2164_),
    .C(_2195_),
    .X(_2426_));
 sky130_fd_sc_hd__a2111o_1 _5793_ (.A1(\mem[12][28] ),
    .A2(_2192_),
    .B1(_2424_),
    .C1(_2425_),
    .D1(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__and3_1 _5794_ (.A(\mem[15][28] ),
    .B(_1494_),
    .C(_2198_),
    .X(_2428_));
 sky130_fd_sc_hd__nor3b_1 _5795_ (.A(_2236_),
    .B(_1601_),
    .C_N(\mem[13][28] ),
    .Y(_2429_));
 sky130_fd_sc_hd__and3_1 _5796_ (.A(\mem[8][28] ),
    .B(_1602_),
    .C(_2170_),
    .X(_2430_));
 sky130_fd_sc_hd__a2111o_1 _5797_ (.A1(\mem[10][28] ),
    .A2(_2234_),
    .B1(_2428_),
    .C1(_2429_),
    .D1(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__nor3_1 _5798_ (.A(_1364_),
    .B(_1607_),
    .C(_1688_),
    .Y(_2432_));
 sky130_fd_sc_hd__and4b_1 _5799_ (.A_N(_1655_),
    .B(_1656_),
    .C(_1610_),
    .D(\mem[22][28] ),
    .X(_2433_));
 sky130_fd_sc_hd__nor3b_1 _5800_ (.A(_2168_),
    .B(_1612_),
    .C_N(\mem[5][28] ),
    .Y(_2434_));
 sky130_fd_sc_hd__a2111o_1 _5801_ (.A1(\mem[1][28] ),
    .A2(_2203_),
    .B1(_2432_),
    .C1(_2433_),
    .D1(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__and3_1 _5802_ (.A(\mem[18][28] ),
    .B(_1504_),
    .C(_1592_),
    .X(_2436_));
 sky130_fd_sc_hd__and3_1 _5803_ (.A(\mem[2][28] ),
    .B(_1616_),
    .C(_1524_),
    .X(_2437_));
 sky130_fd_sc_hd__and3_1 _5804_ (.A(\mem[23][28] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2438_));
 sky130_fd_sc_hd__a2111o_1 _5805_ (.A1(\mem[20][28] ),
    .A2(_2208_),
    .B1(_2436_),
    .C1(_2437_),
    .D1(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__or4_1 _5806_ (.A(_2427_),
    .B(_2431_),
    .C(_2435_),
    .D(_2439_),
    .X(_2440_));
 sky130_fd_sc_hd__a22o_1 _5807_ (.A1(\mem[7][28] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][28] ),
    .X(_2441_));
 sky130_fd_sc_hd__a22o_1 _5808_ (.A1(\mem[31][28] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][28] ),
    .X(_2442_));
 sky130_fd_sc_hd__a22o_1 _5809_ (.A1(\mem[11][28] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][28] ),
    .X(_2443_));
 sky130_fd_sc_hd__a2111o_1 _5810_ (.A1(\mem[26][28] ),
    .A2(_2249_),
    .B1(_2441_),
    .C1(_2442_),
    .D1(_2443_),
    .X(_2444_));
 sky130_fd_sc_hd__a22o_1 _5811_ (.A1(\mem[16][28] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][28] ),
    .X(_2445_));
 sky130_fd_sc_hd__a221o_1 _5812_ (.A1(\mem[6][28] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][28] ),
    .C1(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__a22o_1 _5813_ (.A1(\mem[28][28] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][28] ),
    .X(_2447_));
 sky130_fd_sc_hd__a221o_1 _5814_ (.A1(\mem[17][28] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][28] ),
    .C1(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__or4_4 _5815_ (.A(_2440_),
    .B(_2444_),
    .C(_2446_),
    .D(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__clkbuf_1 _5816_ (.A(_2449_),
    .X(net70));
 sky130_fd_sc_hd__and3_1 _5817_ (.A(\mem[24][29] ),
    .B(_1499_),
    .C(_1522_),
    .X(_2450_));
 sky130_fd_sc_hd__and3_1 _5818_ (.A(\mem[30][29] ),
    .B(_1509_),
    .C(_2174_),
    .X(_2451_));
 sky130_fd_sc_hd__and3_1 _5819_ (.A(\mem[27][29] ),
    .B(_1589_),
    .C(_2195_),
    .X(_2452_));
 sky130_fd_sc_hd__a2111o_1 _5820_ (.A1(\mem[12][29] ),
    .A2(_2192_),
    .B1(_2450_),
    .C1(_2451_),
    .D1(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__and3_1 _5821_ (.A(\mem[15][29] ),
    .B(_1494_),
    .C(_2198_),
    .X(_2454_));
 sky130_fd_sc_hd__nor3b_1 _5822_ (.A(_2236_),
    .B(_1601_),
    .C_N(\mem[13][29] ),
    .Y(_2455_));
 sky130_fd_sc_hd__and3_1 _5823_ (.A(\mem[8][29] ),
    .B(_1602_),
    .C(_1590_),
    .X(_2456_));
 sky130_fd_sc_hd__a2111o_1 _5824_ (.A1(\mem[10][29] ),
    .A2(_2234_),
    .B1(_2454_),
    .C1(_2455_),
    .D1(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__nor3_1 _5825_ (.A(_1399_),
    .B(_1579_),
    .C(_1688_),
    .Y(_2458_));
 sky130_fd_sc_hd__and4b_1 _5826_ (.A_N(_1655_),
    .B(_1656_),
    .C(_1610_),
    .D(\mem[22][29] ),
    .X(_2459_));
 sky130_fd_sc_hd__nor3b_1 _5827_ (.A(_2168_),
    .B(_1612_),
    .C_N(\mem[5][29] ),
    .Y(_2460_));
 sky130_fd_sc_hd__a2111o_1 _5828_ (.A1(\mem[1][29] ),
    .A2(_2203_),
    .B1(_2458_),
    .C1(_2459_),
    .D1(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__and3_1 _5829_ (.A(\mem[18][29] ),
    .B(_1504_),
    .C(_1592_),
    .X(_2462_));
 sky130_fd_sc_hd__and3_1 _5830_ (.A(\mem[2][29] ),
    .B(_1616_),
    .C(_1524_),
    .X(_2463_));
 sky130_fd_sc_hd__and3_1 _5831_ (.A(\mem[23][29] ),
    .B(_2211_),
    .C(_2212_),
    .X(_2464_));
 sky130_fd_sc_hd__a2111o_1 _5832_ (.A1(\mem[20][29] ),
    .A2(_2208_),
    .B1(_2462_),
    .C1(_2463_),
    .D1(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__or4_1 _5833_ (.A(_2453_),
    .B(_2457_),
    .C(_2461_),
    .D(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__a22o_1 _5834_ (.A1(\mem[7][29] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(\mem[9][29] ),
    .X(_2467_));
 sky130_fd_sc_hd__a22o_1 _5835_ (.A1(\mem[31][29] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][29] ),
    .X(_2468_));
 sky130_fd_sc_hd__a22o_1 _5836_ (.A1(\mem[11][29] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][29] ),
    .X(_2469_));
 sky130_fd_sc_hd__a2111o_1 _5837_ (.A1(\mem[26][29] ),
    .A2(_2249_),
    .B1(_2467_),
    .C1(_2468_),
    .D1(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__a22o_1 _5838_ (.A1(\mem[16][29] ),
    .A2(_2222_),
    .B1(_2223_),
    .B2(\mem[19][29] ),
    .X(_2471_));
 sky130_fd_sc_hd__a221o_1 _5839_ (.A1(\mem[6][29] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][29] ),
    .C1(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__a22o_1 _5840_ (.A1(\mem[28][29] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][29] ),
    .X(_2473_));
 sky130_fd_sc_hd__a221o_1 _5841_ (.A1(\mem[17][29] ),
    .A2(_2226_),
    .B1(_2262_),
    .B2(\mem[21][29] ),
    .C1(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__or4_2 _5842_ (.A(_2466_),
    .B(_2470_),
    .C(_2472_),
    .D(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__clkbuf_4 _5843_ (.A(_2475_),
    .X(net71));
 sky130_fd_sc_hd__and3_1 _5844_ (.A(\mem[24][30] ),
    .B(_1499_),
    .C(_1522_),
    .X(_2476_));
 sky130_fd_sc_hd__and3_1 _5845_ (.A(\mem[30][30] ),
    .B(_1509_),
    .C(_2174_),
    .X(_2477_));
 sky130_fd_sc_hd__and3_1 _5846_ (.A(\mem[27][30] ),
    .B(_1589_),
    .C(_1497_),
    .X(_2478_));
 sky130_fd_sc_hd__a2111o_1 _5847_ (.A1(\mem[12][30] ),
    .A2(_1511_),
    .B1(_2476_),
    .C1(_2477_),
    .D1(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__and3_1 _5848_ (.A(\mem[15][30] ),
    .B(_1494_),
    .C(_1500_),
    .X(_2480_));
 sky130_fd_sc_hd__nor3b_1 _5849_ (.A(_2236_),
    .B(_1601_),
    .C_N(\mem[13][30] ),
    .Y(_2481_));
 sky130_fd_sc_hd__and3_1 _5850_ (.A(\mem[8][30] ),
    .B(_1602_),
    .C(_1590_),
    .X(_2482_));
 sky130_fd_sc_hd__a2111o_1 _5851_ (.A1(\mem[10][30] ),
    .A2(_2234_),
    .B1(_2480_),
    .C1(_2481_),
    .D1(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__nor3_1 _5852_ (.A(_1440_),
    .B(_1579_),
    .C(_1549_),
    .Y(_2484_));
 sky130_fd_sc_hd__and4b_1 _5853_ (.A_N(_1655_),
    .B(_1656_),
    .C(_1610_),
    .D(\mem[22][30] ),
    .X(_2485_));
 sky130_fd_sc_hd__nor3b_1 _5854_ (.A(_2168_),
    .B(_1612_),
    .C_N(\mem[5][30] ),
    .Y(_2486_));
 sky130_fd_sc_hd__a2111o_1 _5855_ (.A1(\mem[1][30] ),
    .A2(_1550_),
    .B1(_2484_),
    .C1(_2485_),
    .D1(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__and3_1 _5856_ (.A(\mem[18][30] ),
    .B(_1504_),
    .C(_1592_),
    .X(_2488_));
 sky130_fd_sc_hd__and3_1 _5857_ (.A(\mem[2][30] ),
    .B(_1616_),
    .C(_1524_),
    .X(_2489_));
 sky130_fd_sc_hd__and3_1 _5858_ (.A(\mem[23][30] ),
    .B(_1594_),
    .C(_1564_),
    .X(_2490_));
 sky130_fd_sc_hd__a2111o_1 _5859_ (.A1(\mem[20][30] ),
    .A2(_1541_),
    .B1(_2488_),
    .C1(_2489_),
    .D1(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__or4_1 _5860_ (.A(_2479_),
    .B(_2483_),
    .C(_2487_),
    .D(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__a22o_1 _5861_ (.A1(\mem[7][30] ),
    .A2(_1565_),
    .B1(_1571_),
    .B2(\mem[9][30] ),
    .X(_2493_));
 sky130_fd_sc_hd__a22o_1 _5862_ (.A1(\mem[31][30] ),
    .A2(_2251_),
    .B1(_2252_),
    .B2(\mem[25][30] ),
    .X(_2494_));
 sky130_fd_sc_hd__a22o_1 _5863_ (.A1(\mem[11][30] ),
    .A2(_2254_),
    .B1(_2255_),
    .B2(\mem[14][30] ),
    .X(_2495_));
 sky130_fd_sc_hd__a2111o_1 _5864_ (.A1(\mem[26][30] ),
    .A2(_2249_),
    .B1(_2493_),
    .C1(_2494_),
    .D1(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__a22o_1 _5865_ (.A1(\mem[16][30] ),
    .A2(_1546_),
    .B1(_1580_),
    .B2(\mem[19][30] ),
    .X(_2497_));
 sky130_fd_sc_hd__a221o_1 _5866_ (.A1(\mem[6][30] ),
    .A2(_2258_),
    .B1(_2259_),
    .B2(\mem[4][30] ),
    .C1(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a22o_1 _5867_ (.A1(\mem[28][30] ),
    .A2(_2263_),
    .B1(_2264_),
    .B2(\mem[29][30] ),
    .X(_2499_));
 sky130_fd_sc_hd__a221o_1 _5868_ (.A1(\mem[17][30] ),
    .A2(_1530_),
    .B1(_2262_),
    .B2(\mem[21][30] ),
    .C1(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__or4_4 _5869_ (.A(_2492_),
    .B(_2496_),
    .C(_2498_),
    .D(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__clkbuf_4 _5870_ (.A(_2501_),
    .X(net73));
 sky130_fd_sc_hd__and3_1 _5871_ (.A(\mem[24][31] ),
    .B(_1499_),
    .C(_1522_),
    .X(_2502_));
 sky130_fd_sc_hd__and3_1 _5872_ (.A(\mem[30][31] ),
    .B(_1509_),
    .C(_2174_),
    .X(_2503_));
 sky130_fd_sc_hd__and3_1 _5873_ (.A(\mem[27][31] ),
    .B(_1589_),
    .C(_1497_),
    .X(_2504_));
 sky130_fd_sc_hd__a2111o_1 _5874_ (.A1(\mem[12][31] ),
    .A2(_1511_),
    .B1(_2502_),
    .C1(_2503_),
    .D1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__and3_1 _5875_ (.A(\mem[15][31] ),
    .B(_1494_),
    .C(_1500_),
    .X(_2506_));
 sky130_fd_sc_hd__nor3b_1 _5876_ (.A(_1619_),
    .B(_1601_),
    .C_N(\mem[13][31] ),
    .Y(_2507_));
 sky130_fd_sc_hd__and3_1 _5877_ (.A(\mem[8][31] ),
    .B(_1602_),
    .C(_1590_),
    .X(_2508_));
 sky130_fd_sc_hd__a2111o_1 _5878_ (.A1(\mem[10][31] ),
    .A2(_1597_),
    .B1(_2506_),
    .C1(_2507_),
    .D1(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__and4b_1 _5879_ (.A_N(_1517_),
    .B(_1516_),
    .C(_1657_),
    .D(\mem[22][31] ),
    .X(_2510_));
 sky130_fd_sc_hd__nor3_1 _5880_ (.A(_1473_),
    .B(_2026_),
    .C(_1608_),
    .Y(_2511_));
 sky130_fd_sc_hd__nor3b_1 _5881_ (.A(_2168_),
    .B(_1612_),
    .C_N(\mem[5][31] ),
    .Y(_2512_));
 sky130_fd_sc_hd__a2111o_1 _5882_ (.A1(\mem[1][31] ),
    .A2(_1550_),
    .B1(_2510_),
    .C1(_2511_),
    .D1(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__and3_1 _5883_ (.A(\mem[18][31] ),
    .B(_1504_),
    .C(_1592_),
    .X(_2514_));
 sky130_fd_sc_hd__and3_1 _5884_ (.A(\mem[2][31] ),
    .B(_1616_),
    .C(_1524_),
    .X(_2515_));
 sky130_fd_sc_hd__and3_1 _5885_ (.A(\mem[23][31] ),
    .B(_1594_),
    .C(_1564_),
    .X(_2516_));
 sky130_fd_sc_hd__a2111o_1 _5886_ (.A1(\mem[20][31] ),
    .A2(_1541_),
    .B1(_2514_),
    .C1(_2515_),
    .D1(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__or4_1 _5887_ (.A(_2505_),
    .B(_2509_),
    .C(_2513_),
    .D(_2517_),
    .X(_2518_));
 sky130_fd_sc_hd__a22o_1 _5888_ (.A1(\mem[7][31] ),
    .A2(_1565_),
    .B1(_1571_),
    .B2(\mem[9][31] ),
    .X(_2519_));
 sky130_fd_sc_hd__a22o_1 _5889_ (.A1(\mem[31][31] ),
    .A2(_1501_),
    .B1(_1520_),
    .B2(\mem[25][31] ),
    .X(_2520_));
 sky130_fd_sc_hd__a22o_1 _5890_ (.A1(\mem[11][31] ),
    .A2(_1498_),
    .B1(_1525_),
    .B2(\mem[14][31] ),
    .X(_2521_));
 sky130_fd_sc_hd__a2111o_1 _5891_ (.A1(\mem[26][31] ),
    .A2(_1623_),
    .B1(_2519_),
    .C1(_2520_),
    .D1(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__a22o_1 _5892_ (.A1(\mem[16][31] ),
    .A2(_1546_),
    .B1(_1580_),
    .B2(\mem[19][31] ),
    .X(_2523_));
 sky130_fd_sc_hd__a221o_1 _5893_ (.A1(\mem[6][31] ),
    .A2(_1539_),
    .B1(_1554_),
    .B2(\mem[4][31] ),
    .C1(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__a22o_1 _5894_ (.A1(\mem[28][31] ),
    .A2(_1639_),
    .B1(_1641_),
    .B2(\mem[29][31] ),
    .X(_2525_));
 sky130_fd_sc_hd__a221o_1 _5895_ (.A1(\mem[17][31] ),
    .A2(_1530_),
    .B1(_1637_),
    .B2(\mem[21][31] ),
    .C1(_2525_),
    .X(_2526_));
 sky130_fd_sc_hd__or4_4 _5896_ (.A(_2518_),
    .B(_2522_),
    .C(_2524_),
    .D(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__clkbuf_1 _5897_ (.A(_2527_),
    .X(net74));
 sky130_fd_sc_hd__and3_1 _5898_ (.A(\mem[6][0] ),
    .B(_1044_),
    .C(_1058_),
    .X(_2528_));
 sky130_fd_sc_hd__and3_1 _5899_ (.A(\mem[28][0] ),
    .B(_1001_),
    .C(_1062_),
    .X(_2529_));
 sky130_fd_sc_hd__and3_1 _5900_ (.A(\mem[4][0] ),
    .B(_1052_),
    .C(_1055_),
    .X(_2530_));
 sky130_fd_sc_hd__a2111o_1 _5901_ (.A1(\mem[2][0] ),
    .A2(_1092_),
    .B1(_2528_),
    .C1(_2529_),
    .D1(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__and3_1 _5902_ (.A(\mem[31][0] ),
    .B(_1067_),
    .C(_1235_),
    .X(_2532_));
 sky130_fd_sc_hd__nor3b_1 _5903_ (.A(_1073_),
    .B(_1041_),
    .C_N(\mem[5][0] ),
    .Y(_2533_));
 sky130_fd_sc_hd__and3_1 _5904_ (.A(\mem[29][0] ),
    .B(_1011_),
    .C(_1396_),
    .X(_2534_));
 sky130_fd_sc_hd__a2111o_1 _5905_ (.A1(\mem[26][0] ),
    .A2(_1068_),
    .B1(_2532_),
    .C1(_2533_),
    .D1(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__nor3_1 _5906_ (.A(_1555_),
    .B(_1045_),
    .C(_1041_),
    .Y(_2536_));
 sky130_fd_sc_hd__and3_1 _5907_ (.A(\mem[12][0] ),
    .B(_1001_),
    .C(_1004_),
    .X(_2537_));
 sky130_fd_sc_hd__inv_2 _5908_ (.A(\mem[19][0] ),
    .Y(_2538_));
 sky130_fd_sc_hd__nor3_1 _5909_ (.A(_2538_),
    .B(_1045_),
    .C(_1046_),
    .Y(_2539_));
 sky130_fd_sc_hd__a2111o_1 _5910_ (.A1(\mem[17][0] ),
    .A2(_1098_),
    .B1(_2536_),
    .C1(_2537_),
    .D1(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__and3_1 _5911_ (.A(\mem[20][0] ),
    .B(_1055_),
    .C(_1024_),
    .X(_2541_));
 sky130_fd_sc_hd__and3_1 _5912_ (.A(\mem[15][0] ),
    .B(_1026_),
    .C(_1028_),
    .X(_2542_));
 sky130_fd_sc_hd__and3_1 _5913_ (.A(\mem[13][0] ),
    .B(_1026_),
    .C(_1110_),
    .X(_2543_));
 sky130_fd_sc_hd__a2111o_1 _5914_ (.A1(\mem[11][0] ),
    .A2(_1078_),
    .B1(_2541_),
    .C1(_2542_),
    .D1(_2543_),
    .X(_2544_));
 sky130_fd_sc_hd__or4_1 _5915_ (.A(_2531_),
    .B(_2535_),
    .C(_2540_),
    .D(_2544_),
    .X(_2545_));
 sky130_fd_sc_hd__a22o_1 _5916_ (.A1(\mem[25][0] ),
    .A2(_0997_),
    .B1(_1128_),
    .B2(\mem[27][0] ),
    .X(_2546_));
 sky130_fd_sc_hd__nor2_1 _5917_ (.A(_1073_),
    .B(_1046_),
    .Y(_2547_));
 sky130_fd_sc_hd__a22o_1 _5918_ (.A1(\mem[8][0] ),
    .A2(_1082_),
    .B1(_2547_),
    .B2(\mem[3][0] ),
    .X(_2548_));
 sky130_fd_sc_hd__nor2_1 _5919_ (.A(_1073_),
    .B(_1119_),
    .Y(_2549_));
 sky130_fd_sc_hd__a32o_1 _5920_ (.A1(\mem[30][0] ),
    .A2(_1073_),
    .A3(_1013_),
    .B1(_2549_),
    .B2(\mem[1][0] ),
    .X(_2550_));
 sky130_fd_sc_hd__a2111o_1 _5921_ (.A1(\mem[7][0] ),
    .A2(_1089_),
    .B1(_2546_),
    .C1(_2548_),
    .D1(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__and3_1 _5922_ (.A(\mem[22][0] ),
    .B(_1073_),
    .C(_1059_),
    .X(_2552_));
 sky130_fd_sc_hd__a31o_1 _5923_ (.A1(\mem[24][0] ),
    .A2(_1022_),
    .A3(_1063_),
    .B1(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a221o_1 _5924_ (.A1(\mem[9][0] ),
    .A2(_1077_),
    .B1(_1094_),
    .B2(\mem[23][0] ),
    .C1(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__a22o_1 _5925_ (.A1(\mem[14][0] ),
    .A2(_1133_),
    .B1(_1017_),
    .B2(\mem[10][0] ),
    .X(_2555_));
 sky130_fd_sc_hd__a221o_1 _5926_ (.A1(\mem[18][0] ),
    .A2(_1051_),
    .B1(_1087_),
    .B2(\mem[16][0] ),
    .C1(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__or4_4 _5927_ (.A(_2545_),
    .B(_2551_),
    .C(_2554_),
    .D(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__clkbuf_1 _5928_ (.A(_2557_),
    .X(net82));
 sky130_fd_sc_hd__and3_1 _5929_ (.A(\mem[12][1] ),
    .B(_1319_),
    .C(_1260_),
    .X(_2558_));
 sky130_fd_sc_hd__and3_1 _5930_ (.A(\mem[29][1] ),
    .B(_1202_),
    .C(_1321_),
    .X(_2559_));
 sky130_fd_sc_hd__and3_1 _5931_ (.A(\mem[30][1] ),
    .B(_1232_),
    .C(_1356_),
    .X(_2560_));
 sky130_fd_sc_hd__a2111o_1 _5932_ (.A1(\mem[25][1] ),
    .A2(_1353_),
    .B1(_2558_),
    .C1(_2559_),
    .D1(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__and3_1 _5933_ (.A(\mem[15][1] ),
    .B(_1435_),
    .C(_1235_),
    .X(_2562_));
 sky130_fd_sc_hd__and3_1 _5934_ (.A(\mem[24][1] ),
    .B(_1326_),
    .C(_1295_),
    .X(_2563_));
 sky130_fd_sc_hd__and3_1 _5935_ (.A(\mem[13][1] ),
    .B(_1470_),
    .C(_1396_),
    .X(_2564_));
 sky130_fd_sc_hd__a2111o_1 _5936_ (.A1(\mem[10][1] ),
    .A2(_1359_),
    .B1(_2562_),
    .C1(_2563_),
    .D1(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__inv_2 _5937_ (.A(\mem[19][1] ),
    .Y(_2566_));
 sky130_fd_sc_hd__or3_1 _5938_ (.A(_2566_),
    .B(_1115_),
    .C(_1152_),
    .X(_2567_));
 sky130_fd_sc_hd__buf_2 _5939_ (.A(_1010_),
    .X(_2568_));
 sky130_fd_sc_hd__or3b_1 _5940_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][1] ),
    .X(_2569_));
 sky130_fd_sc_hd__or3b_1 _5941_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][1] ),
    .X(_2570_));
 sky130_fd_sc_hd__o2111ai_1 _5942_ (.A1(_1606_),
    .A2(_1400_),
    .B1(_2567_),
    .C1(_2569_),
    .D1(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__and3_1 _5943_ (.A(\mem[4][1] ),
    .B(_1336_),
    .C(_1275_),
    .X(_2572_));
 sky130_fd_sc_hd__and3_1 _5944_ (.A(\mem[22][1] ),
    .B(_1338_),
    .C(_1339_),
    .X(_2573_));
 sky130_fd_sc_hd__and3_1 _5945_ (.A(\mem[20][1] ),
    .B(_1373_),
    .C(_1374_),
    .X(_2574_));
 sky130_fd_sc_hd__a2111o_1 _5946_ (.A1(\mem[18][1] ),
    .A2(_1370_),
    .B1(_2572_),
    .C1(_2573_),
    .D1(_2574_),
    .X(_2575_));
 sky130_fd_sc_hd__or4_1 _5947_ (.A(_2561_),
    .B(_2565_),
    .C(_2571_),
    .D(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__a22o_1 _5948_ (.A1(\mem[9][1] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][1] ),
    .X(_2577_));
 sky130_fd_sc_hd__a22o_1 _5949_ (.A1(\mem[27][1] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][1] ),
    .X(_2578_));
 sky130_fd_sc_hd__buf_6 _5950_ (.A(_1073_),
    .X(_2579_));
 sky130_fd_sc_hd__a32o_1 _5951_ (.A1(_2579_),
    .A2(\mem[31][1] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][1] ),
    .X(_2580_));
 sky130_fd_sc_hd__a2111o_1 _5952_ (.A1(\mem[26][1] ),
    .A2(_1412_),
    .B1(_2577_),
    .C1(_2578_),
    .D1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__a22o_1 _5953_ (.A1(\mem[16][1] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][1] ),
    .X(_2582_));
 sky130_fd_sc_hd__a221o_1 _5954_ (.A1(\mem[8][1] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][1] ),
    .C1(_2582_),
    .X(_2583_));
 sky130_fd_sc_hd__a22o_1 _5955_ (.A1(\mem[21][1] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][1] ),
    .X(_2584_));
 sky130_fd_sc_hd__a221o_1 _5956_ (.A1(\mem[2][1] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][1] ),
    .C1(_2584_),
    .X(_2585_));
 sky130_fd_sc_hd__or4_4 _5957_ (.A(_2576_),
    .B(_2581_),
    .C(_2583_),
    .D(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _5958_ (.A(_2586_),
    .X(net93));
 sky130_fd_sc_hd__and3_1 _5959_ (.A(\mem[12][2] ),
    .B(_1319_),
    .C(_1260_),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_4 _5960_ (.A(_0995_),
    .X(_2588_));
 sky130_fd_sc_hd__and3_1 _5961_ (.A(\mem[29][2] ),
    .B(_2588_),
    .C(_1321_),
    .X(_2589_));
 sky130_fd_sc_hd__and3_1 _5962_ (.A(\mem[30][2] ),
    .B(_1232_),
    .C(_1356_),
    .X(_2590_));
 sky130_fd_sc_hd__a2111o_1 _5963_ (.A1(\mem[25][2] ),
    .A2(_1353_),
    .B1(_2587_),
    .C1(_2589_),
    .D1(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_4 _5964_ (.A(_1027_),
    .X(_2592_));
 sky130_fd_sc_hd__and3_1 _5965_ (.A(\mem[15][2] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2593_));
 sky130_fd_sc_hd__and3_1 _5966_ (.A(\mem[24][2] ),
    .B(_1326_),
    .C(_1295_),
    .X(_2594_));
 sky130_fd_sc_hd__and3_1 _5967_ (.A(\mem[13][2] ),
    .B(_1470_),
    .C(_1396_),
    .X(_2595_));
 sky130_fd_sc_hd__a2111o_1 _5968_ (.A1(\mem[10][2] ),
    .A2(_1359_),
    .B1(_2593_),
    .C1(_2594_),
    .D1(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__inv_2 _5969_ (.A(\mem[19][2] ),
    .Y(_2597_));
 sky130_fd_sc_hd__clkbuf_4 _5970_ (.A(_1044_),
    .X(_2598_));
 sky130_fd_sc_hd__or3_1 _5971_ (.A(_2597_),
    .B(_2598_),
    .C(_1152_),
    .X(_2599_));
 sky130_fd_sc_hd__or3b_1 _5972_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][2] ),
    .X(_2600_));
 sky130_fd_sc_hd__or3b_1 _5973_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][2] ),
    .X(_2601_));
 sky130_fd_sc_hd__o2111ai_2 _5974_ (.A1(_1659_),
    .A2(_1400_),
    .B1(_2599_),
    .C1(_2600_),
    .D1(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__and3_1 _5975_ (.A(\mem[4][2] ),
    .B(_1336_),
    .C(_1275_),
    .X(_2603_));
 sky130_fd_sc_hd__and3_1 _5976_ (.A(\mem[22][2] ),
    .B(_1338_),
    .C(_1339_),
    .X(_2604_));
 sky130_fd_sc_hd__and3_1 _5977_ (.A(\mem[20][2] ),
    .B(_1373_),
    .C(_1374_),
    .X(_2605_));
 sky130_fd_sc_hd__a2111o_1 _5978_ (.A1(\mem[18][2] ),
    .A2(_1370_),
    .B1(_2603_),
    .C1(_2604_),
    .D1(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__or4_1 _5979_ (.A(_2591_),
    .B(_2596_),
    .C(_2602_),
    .D(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__a22o_1 _5980_ (.A1(\mem[9][2] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][2] ),
    .X(_2608_));
 sky130_fd_sc_hd__a22o_1 _5981_ (.A1(\mem[27][2] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][2] ),
    .X(_2609_));
 sky130_fd_sc_hd__a32o_1 _5982_ (.A1(_2579_),
    .A2(\mem[31][2] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][2] ),
    .X(_2610_));
 sky130_fd_sc_hd__a2111o_1 _5983_ (.A1(\mem[26][2] ),
    .A2(_1412_),
    .B1(_2608_),
    .C1(_2609_),
    .D1(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__a22o_1 _5984_ (.A1(\mem[16][2] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][2] ),
    .X(_2612_));
 sky130_fd_sc_hd__a221o_1 _5985_ (.A1(\mem[8][2] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][2] ),
    .C1(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__a22o_1 _5986_ (.A1(\mem[21][2] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][2] ),
    .X(_2614_));
 sky130_fd_sc_hd__a221o_1 _5987_ (.A1(\mem[2][2] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][2] ),
    .C1(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__or4_4 _5988_ (.A(_2607_),
    .B(_2611_),
    .C(_2613_),
    .D(_2615_),
    .X(_2616_));
 sky130_fd_sc_hd__buf_4 _5989_ (.A(_2616_),
    .X(net104));
 sky130_fd_sc_hd__and3_1 _5990_ (.A(\mem[12][3] ),
    .B(_1319_),
    .C(_1260_),
    .X(_2617_));
 sky130_fd_sc_hd__and3_1 _5991_ (.A(\mem[29][3] ),
    .B(_2588_),
    .C(_1321_),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_4 _5992_ (.A(_0995_),
    .X(_2619_));
 sky130_fd_sc_hd__and3_1 _5993_ (.A(\mem[30][3] ),
    .B(_2619_),
    .C(_1356_),
    .X(_2620_));
 sky130_fd_sc_hd__a2111o_1 _5994_ (.A1(\mem[25][3] ),
    .A2(_1353_),
    .B1(_2617_),
    .C1(_2618_),
    .D1(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__and3_1 _5995_ (.A(\mem[15][3] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2622_));
 sky130_fd_sc_hd__and3_1 _5996_ (.A(\mem[24][3] ),
    .B(_1326_),
    .C(_1295_),
    .X(_2623_));
 sky130_fd_sc_hd__and3_1 _5997_ (.A(\mem[13][3] ),
    .B(_1470_),
    .C(_1396_),
    .X(_2624_));
 sky130_fd_sc_hd__a2111o_1 _5998_ (.A1(\mem[10][3] ),
    .A2(_1359_),
    .B1(_2622_),
    .C1(_2623_),
    .D1(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__or3b_1 _5999_ (.A(_1036_),
    .B(_1040_),
    .C_N(\mem[5][3] ),
    .X(_2626_));
 sky130_fd_sc_hd__inv_2 _6000_ (.A(\mem[19][3] ),
    .Y(_2627_));
 sky130_fd_sc_hd__or3_1 _6001_ (.A(_2627_),
    .B(_1045_),
    .C(_1046_),
    .X(_2628_));
 sky130_fd_sc_hd__or3b_1 _6002_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][3] ),
    .X(_2629_));
 sky130_fd_sc_hd__o2111ai_2 _6003_ (.A1(_1687_),
    .A2(_1400_),
    .B1(_2626_),
    .C1(_2628_),
    .D1(_2629_),
    .Y(_2630_));
 sky130_fd_sc_hd__and3_1 _6004_ (.A(\mem[4][3] ),
    .B(_1336_),
    .C(_1275_),
    .X(_2631_));
 sky130_fd_sc_hd__and3_1 _6005_ (.A(\mem[22][3] ),
    .B(_1338_),
    .C(_1339_),
    .X(_2632_));
 sky130_fd_sc_hd__and3_1 _6006_ (.A(\mem[20][3] ),
    .B(_1373_),
    .C(_1374_),
    .X(_2633_));
 sky130_fd_sc_hd__a2111o_1 _6007_ (.A1(\mem[18][3] ),
    .A2(_1370_),
    .B1(_2631_),
    .C1(_2632_),
    .D1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__or4_1 _6008_ (.A(_2621_),
    .B(_2625_),
    .C(_2630_),
    .D(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__a22o_1 _6009_ (.A1(\mem[9][3] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][3] ),
    .X(_2636_));
 sky130_fd_sc_hd__a22o_1 _6010_ (.A1(\mem[27][3] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][3] ),
    .X(_2637_));
 sky130_fd_sc_hd__a32o_1 _6011_ (.A1(_2579_),
    .A2(\mem[31][3] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][3] ),
    .X(_2638_));
 sky130_fd_sc_hd__a2111o_1 _6012_ (.A1(\mem[26][3] ),
    .A2(_1412_),
    .B1(_2636_),
    .C1(_2637_),
    .D1(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__a22o_1 _6013_ (.A1(\mem[16][3] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][3] ),
    .X(_2640_));
 sky130_fd_sc_hd__a221o_1 _6014_ (.A1(\mem[8][3] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][3] ),
    .C1(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__a22o_1 _6015_ (.A1(\mem[21][3] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][3] ),
    .X(_2642_));
 sky130_fd_sc_hd__a221o_1 _6016_ (.A1(\mem[2][3] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][3] ),
    .C1(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__or4_4 _6017_ (.A(_2635_),
    .B(_2639_),
    .C(_2641_),
    .D(_2643_),
    .X(_2644_));
 sky130_fd_sc_hd__clkbuf_1 _6018_ (.A(_2644_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 _6019_ (.A(_1002_),
    .X(_2645_));
 sky130_fd_sc_hd__and3_1 _6020_ (.A(\mem[12][4] ),
    .B(_1319_),
    .C(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__and3_1 _6021_ (.A(\mem[29][4] ),
    .B(_2588_),
    .C(_1321_),
    .X(_2647_));
 sky130_fd_sc_hd__and3_1 _6022_ (.A(\mem[30][4] ),
    .B(_2619_),
    .C(_1356_),
    .X(_2648_));
 sky130_fd_sc_hd__a2111o_1 _6023_ (.A1(\mem[25][4] ),
    .A2(_1353_),
    .B1(_2646_),
    .C1(_2647_),
    .D1(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__and3_1 _6024_ (.A(\mem[15][4] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2650_));
 sky130_fd_sc_hd__and3_1 _6025_ (.A(\mem[24][4] ),
    .B(_1326_),
    .C(_1295_),
    .X(_2651_));
 sky130_fd_sc_hd__and3_1 _6026_ (.A(\mem[13][4] ),
    .B(_1470_),
    .C(_1396_),
    .X(_2652_));
 sky130_fd_sc_hd__a2111o_1 _6027_ (.A1(\mem[10][4] ),
    .A2(_1359_),
    .B1(_2650_),
    .C1(_2651_),
    .D1(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__inv_2 _6028_ (.A(\mem[19][4] ),
    .Y(_2654_));
 sky130_fd_sc_hd__buf_2 _6029_ (.A(_1032_),
    .X(_2655_));
 sky130_fd_sc_hd__or3_1 _6030_ (.A(_2654_),
    .B(_2598_),
    .C(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__or3b_1 _6031_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][4] ),
    .X(_2657_));
 sky130_fd_sc_hd__or3b_1 _6032_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][4] ),
    .X(_2658_));
 sky130_fd_sc_hd__o2111ai_2 _6033_ (.A1(_1716_),
    .A2(_1400_),
    .B1(_2656_),
    .C1(_2657_),
    .D1(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__buf_4 _6034_ (.A(_1053_),
    .X(_2660_));
 sky130_fd_sc_hd__and3_1 _6035_ (.A(\mem[4][4] ),
    .B(_1336_),
    .C(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__and3_1 _6036_ (.A(\mem[22][4] ),
    .B(_1338_),
    .C(_1339_),
    .X(_2662_));
 sky130_fd_sc_hd__and3_1 _6037_ (.A(\mem[20][4] ),
    .B(_1373_),
    .C(_1374_),
    .X(_2663_));
 sky130_fd_sc_hd__a2111o_1 _6038_ (.A1(\mem[18][4] ),
    .A2(_1370_),
    .B1(_2661_),
    .C1(_2662_),
    .D1(_2663_),
    .X(_2664_));
 sky130_fd_sc_hd__or4_1 _6039_ (.A(_2649_),
    .B(_2653_),
    .C(_2659_),
    .D(_2664_),
    .X(_2665_));
 sky130_fd_sc_hd__a22o_1 _6040_ (.A1(\mem[9][4] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][4] ),
    .X(_2666_));
 sky130_fd_sc_hd__a22o_1 _6041_ (.A1(\mem[27][4] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][4] ),
    .X(_2667_));
 sky130_fd_sc_hd__a32o_1 _6042_ (.A1(_2579_),
    .A2(\mem[31][4] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][4] ),
    .X(_2668_));
 sky130_fd_sc_hd__a2111o_1 _6043_ (.A1(\mem[26][4] ),
    .A2(_1412_),
    .B1(_2666_),
    .C1(_2667_),
    .D1(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__a22o_1 _6044_ (.A1(\mem[16][4] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][4] ),
    .X(_2670_));
 sky130_fd_sc_hd__a221o_1 _6045_ (.A1(\mem[8][4] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][4] ),
    .C1(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__a22o_1 _6046_ (.A1(\mem[21][4] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][4] ),
    .X(_2672_));
 sky130_fd_sc_hd__a221o_1 _6047_ (.A1(\mem[2][4] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][4] ),
    .C1(_2672_),
    .X(_2673_));
 sky130_fd_sc_hd__or4_4 _6048_ (.A(_2665_),
    .B(_2669_),
    .C(_2671_),
    .D(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__clkbuf_1 _6049_ (.A(_2674_),
    .X(net108));
 sky130_fd_sc_hd__and3_1 _6050_ (.A(\mem[12][5] ),
    .B(_1319_),
    .C(_2645_),
    .X(_2675_));
 sky130_fd_sc_hd__and3_1 _6051_ (.A(\mem[29][5] ),
    .B(_2588_),
    .C(_1321_),
    .X(_2676_));
 sky130_fd_sc_hd__and3_1 _6052_ (.A(\mem[30][5] ),
    .B(_2619_),
    .C(_1356_),
    .X(_2677_));
 sky130_fd_sc_hd__a2111o_1 _6053_ (.A1(\mem[25][5] ),
    .A2(_1353_),
    .B1(_2675_),
    .C1(_2676_),
    .D1(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__and3_1 _6054_ (.A(\mem[15][5] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2679_));
 sky130_fd_sc_hd__clkbuf_4 _6055_ (.A(_1023_),
    .X(_2680_));
 sky130_fd_sc_hd__and3_1 _6056_ (.A(\mem[24][5] ),
    .B(_1326_),
    .C(_2680_),
    .X(_2681_));
 sky130_fd_sc_hd__and3_1 _6057_ (.A(\mem[13][5] ),
    .B(_1470_),
    .C(_1396_),
    .X(_2682_));
 sky130_fd_sc_hd__a2111o_1 _6058_ (.A1(\mem[10][5] ),
    .A2(_1359_),
    .B1(_2679_),
    .C1(_2681_),
    .D1(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__inv_2 _6059_ (.A(\mem[19][5] ),
    .Y(_2684_));
 sky130_fd_sc_hd__or3_1 _6060_ (.A(_2684_),
    .B(_2598_),
    .C(_2655_),
    .X(_2685_));
 sky130_fd_sc_hd__or3b_1 _6061_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][5] ),
    .X(_2686_));
 sky130_fd_sc_hd__or3b_1 _6062_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][5] ),
    .X(_2687_));
 sky130_fd_sc_hd__o2111ai_1 _6063_ (.A1(_1747_),
    .A2(_1400_),
    .B1(_2685_),
    .C1(_2686_),
    .D1(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__and3_1 _6064_ (.A(\mem[4][5] ),
    .B(_1336_),
    .C(_2660_),
    .X(_2689_));
 sky130_fd_sc_hd__and3_1 _6065_ (.A(\mem[22][5] ),
    .B(_1338_),
    .C(_1339_),
    .X(_2690_));
 sky130_fd_sc_hd__and3_1 _6066_ (.A(\mem[20][5] ),
    .B(_1373_),
    .C(_1374_),
    .X(_2691_));
 sky130_fd_sc_hd__a2111o_1 _6067_ (.A1(\mem[18][5] ),
    .A2(_1370_),
    .B1(_2689_),
    .C1(_2690_),
    .D1(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__or4_1 _6068_ (.A(_2678_),
    .B(_2683_),
    .C(_2688_),
    .D(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__a22o_1 _6069_ (.A1(\mem[9][5] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][5] ),
    .X(_2694_));
 sky130_fd_sc_hd__a22o_1 _6070_ (.A1(\mem[27][5] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][5] ),
    .X(_2695_));
 sky130_fd_sc_hd__a32o_1 _6071_ (.A1(_2579_),
    .A2(\mem[31][5] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][5] ),
    .X(_2696_));
 sky130_fd_sc_hd__a2111o_1 _6072_ (.A1(\mem[26][5] ),
    .A2(_1412_),
    .B1(_2694_),
    .C1(_2695_),
    .D1(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__a22o_1 _6073_ (.A1(\mem[16][5] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][5] ),
    .X(_2698_));
 sky130_fd_sc_hd__a221o_1 _6074_ (.A1(\mem[8][5] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][5] ),
    .C1(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__a22o_1 _6075_ (.A1(\mem[21][5] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][5] ),
    .X(_2700_));
 sky130_fd_sc_hd__a221o_1 _6076_ (.A1(\mem[2][5] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][5] ),
    .C1(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__or4_4 _6077_ (.A(_2693_),
    .B(_2697_),
    .C(_2699_),
    .D(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__clkbuf_1 _6078_ (.A(_2702_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 _6079_ (.A(_1000_),
    .X(_2703_));
 sky130_fd_sc_hd__and3_1 _6080_ (.A(\mem[12][6] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2704_));
 sky130_fd_sc_hd__clkbuf_4 _6081_ (.A(_1007_),
    .X(_2705_));
 sky130_fd_sc_hd__and3_1 _6082_ (.A(\mem[29][6] ),
    .B(_2588_),
    .C(_2705_),
    .X(_2706_));
 sky130_fd_sc_hd__and3_1 _6083_ (.A(\mem[30][6] ),
    .B(_2619_),
    .C(_1356_),
    .X(_2707_));
 sky130_fd_sc_hd__a2111o_1 _6084_ (.A1(\mem[25][6] ),
    .A2(_1353_),
    .B1(_2704_),
    .C1(_2706_),
    .D1(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__and3_1 _6085_ (.A(\mem[15][6] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2709_));
 sky130_fd_sc_hd__clkbuf_4 _6086_ (.A(_1021_),
    .X(_2710_));
 sky130_fd_sc_hd__and3_1 _6087_ (.A(\mem[24][6] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2711_));
 sky130_fd_sc_hd__and3_1 _6088_ (.A(\mem[13][6] ),
    .B(_1470_),
    .C(_1396_),
    .X(_2712_));
 sky130_fd_sc_hd__a2111o_1 _6089_ (.A1(\mem[10][6] ),
    .A2(_1359_),
    .B1(_2709_),
    .C1(_2711_),
    .D1(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__or3b_1 _6090_ (.A(_1057_),
    .B(_1040_),
    .C_N(\mem[5][6] ),
    .X(_2714_));
 sky130_fd_sc_hd__inv_2 _6091_ (.A(\mem[19][6] ),
    .Y(_2715_));
 sky130_fd_sc_hd__or3_1 _6092_ (.A(_2715_),
    .B(_1045_),
    .C(_1046_),
    .X(_2716_));
 sky130_fd_sc_hd__or3b_1 _6093_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][6] ),
    .X(_2717_));
 sky130_fd_sc_hd__o2111ai_1 _6094_ (.A1(_1775_),
    .A2(_1400_),
    .B1(_2714_),
    .C1(_2716_),
    .D1(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__clkbuf_4 _6095_ (.A(_1003_),
    .X(_2719_));
 sky130_fd_sc_hd__and3_1 _6096_ (.A(\mem[4][6] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2720_));
 sky130_fd_sc_hd__clkbuf_4 _6097_ (.A(_0995_),
    .X(_2721_));
 sky130_fd_sc_hd__clkbuf_4 _6098_ (.A(_1058_),
    .X(_2722_));
 sky130_fd_sc_hd__and3_1 _6099_ (.A(\mem[22][6] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__and3_1 _6100_ (.A(\mem[20][6] ),
    .B(_1373_),
    .C(_1374_),
    .X(_2724_));
 sky130_fd_sc_hd__a2111o_1 _6101_ (.A1(\mem[18][6] ),
    .A2(_1370_),
    .B1(_2720_),
    .C1(_2723_),
    .D1(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__or4_1 _6102_ (.A(_2708_),
    .B(_2713_),
    .C(_2718_),
    .D(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__a22o_1 _6103_ (.A1(\mem[9][6] ),
    .A2(_1378_),
    .B1(_1413_),
    .B2(\mem[11][6] ),
    .X(_2727_));
 sky130_fd_sc_hd__a22o_1 _6104_ (.A1(\mem[27][6] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][6] ),
    .X(_2728_));
 sky130_fd_sc_hd__a32o_1 _6105_ (.A1(_2579_),
    .A2(\mem[31][6] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][6] ),
    .X(_2729_));
 sky130_fd_sc_hd__a2111o_1 _6106_ (.A1(\mem[26][6] ),
    .A2(_1412_),
    .B1(_2727_),
    .C1(_2728_),
    .D1(_2729_),
    .X(_2730_));
 sky130_fd_sc_hd__a22o_1 _6107_ (.A1(\mem[16][6] ),
    .A2(_1383_),
    .B1(_1384_),
    .B2(\mem[7][6] ),
    .X(_2731_));
 sky130_fd_sc_hd__a221o_1 _6108_ (.A1(\mem[8][6] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][6] ),
    .C1(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__a22o_1 _6109_ (.A1(\mem[21][6] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][6] ),
    .X(_2733_));
 sky130_fd_sc_hd__a221o_1 _6110_ (.A1(\mem[2][6] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][6] ),
    .C1(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__or4_2 _6111_ (.A(_2726_),
    .B(_2730_),
    .C(_2732_),
    .D(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__buf_2 _6112_ (.A(_2735_),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 _6113_ (.A(_0996_),
    .X(_2736_));
 sky130_fd_sc_hd__and3_1 _6114_ (.A(\mem[12][7] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2737_));
 sky130_fd_sc_hd__and3_1 _6115_ (.A(\mem[29][7] ),
    .B(_2588_),
    .C(_2705_),
    .X(_2738_));
 sky130_fd_sc_hd__clkbuf_4 _6116_ (.A(_1012_),
    .X(_2739_));
 sky130_fd_sc_hd__and3_1 _6117_ (.A(\mem[30][7] ),
    .B(_2619_),
    .C(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__a2111o_1 _6118_ (.A1(\mem[25][7] ),
    .A2(_2736_),
    .B1(_2737_),
    .C1(_2738_),
    .D1(_2740_),
    .X(_2741_));
 sky130_fd_sc_hd__clkbuf_4 _6119_ (.A(_1016_),
    .X(_2742_));
 sky130_fd_sc_hd__and3_1 _6120_ (.A(\mem[15][7] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2743_));
 sky130_fd_sc_hd__and3_1 _6121_ (.A(\mem[24][7] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2744_));
 sky130_fd_sc_hd__buf_2 _6122_ (.A(_1007_),
    .X(_2745_));
 sky130_fd_sc_hd__and3_1 _6123_ (.A(\mem[13][7] ),
    .B(_1470_),
    .C(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__a2111o_1 _6124_ (.A1(\mem[10][7] ),
    .A2(_2742_),
    .B1(_2743_),
    .C1(_2744_),
    .D1(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__inv_2 _6125_ (.A(\mem[19][7] ),
    .Y(_2748_));
 sky130_fd_sc_hd__or3_1 _6126_ (.A(_2748_),
    .B(_2598_),
    .C(_2655_),
    .X(_2749_));
 sky130_fd_sc_hd__or3b_1 _6127_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][7] ),
    .X(_2750_));
 sky130_fd_sc_hd__or3b_1 _6128_ (.A(_1445_),
    .B(_1404_),
    .C_N(\mem[1][7] ),
    .X(_2751_));
 sky130_fd_sc_hd__o2111ai_1 _6129_ (.A1(_1802_),
    .A2(_1400_),
    .B1(_2749_),
    .C1(_2750_),
    .D1(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__clkbuf_4 _6130_ (.A(_1050_),
    .X(_2753_));
 sky130_fd_sc_hd__and3_1 _6131_ (.A(\mem[4][7] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2754_));
 sky130_fd_sc_hd__and3_1 _6132_ (.A(\mem[22][7] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2755_));
 sky130_fd_sc_hd__buf_2 _6133_ (.A(_1054_),
    .X(_2756_));
 sky130_fd_sc_hd__buf_2 _6134_ (.A(_1062_),
    .X(_2757_));
 sky130_fd_sc_hd__and3_1 _6135_ (.A(\mem[20][7] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__a2111o_1 _6136_ (.A1(\mem[18][7] ),
    .A2(_2753_),
    .B1(_2754_),
    .C1(_2755_),
    .D1(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__or4_1 _6137_ (.A(_2741_),
    .B(_2747_),
    .C(_2752_),
    .D(_2759_),
    .X(_2760_));
 sky130_fd_sc_hd__buf_4 _6138_ (.A(_1076_),
    .X(_2761_));
 sky130_fd_sc_hd__a22o_1 _6139_ (.A1(\mem[9][7] ),
    .A2(_2761_),
    .B1(_1413_),
    .B2(\mem[11][7] ),
    .X(_2762_));
 sky130_fd_sc_hd__a22o_1 _6140_ (.A1(\mem[27][7] ),
    .A2(_1415_),
    .B1(_1454_),
    .B2(\mem[28][7] ),
    .X(_2763_));
 sky130_fd_sc_hd__a32o_1 _6141_ (.A1(_2579_),
    .A2(\mem[31][7] ),
    .A3(_1456_),
    .B1(_1417_),
    .B2(\mem[14][7] ),
    .X(_2764_));
 sky130_fd_sc_hd__a2111o_1 _6142_ (.A1(\mem[26][7] ),
    .A2(_1412_),
    .B1(_2762_),
    .C1(_2763_),
    .D1(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__buf_4 _6143_ (.A(_1086_),
    .X(_2766_));
 sky130_fd_sc_hd__buf_4 _6144_ (.A(_1088_),
    .X(_2767_));
 sky130_fd_sc_hd__a22o_1 _6145_ (.A1(\mem[16][7] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][7] ),
    .X(_2768_));
 sky130_fd_sc_hd__a221o_1 _6146_ (.A1(\mem[8][7] ),
    .A2(_1420_),
    .B1(_1421_),
    .B2(\mem[6][7] ),
    .C1(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__a22o_1 _6147_ (.A1(\mem[21][7] ),
    .A2(_1426_),
    .B1(_1427_),
    .B2(\mem[17][7] ),
    .X(_2770_));
 sky130_fd_sc_hd__a221o_1 _6148_ (.A1(\mem[2][7] ),
    .A2(_1424_),
    .B1(_1425_),
    .B2(\mem[23][7] ),
    .C1(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__or4_4 _6149_ (.A(_2760_),
    .B(_2765_),
    .C(_2769_),
    .D(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__buf_4 _6150_ (.A(_2772_),
    .X(net111));
 sky130_fd_sc_hd__and3_1 _6151_ (.A(\mem[12][8] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2773_));
 sky130_fd_sc_hd__and3_1 _6152_ (.A(\mem[29][8] ),
    .B(_2588_),
    .C(_2705_),
    .X(_2774_));
 sky130_fd_sc_hd__and3_1 _6153_ (.A(\mem[30][8] ),
    .B(_2619_),
    .C(_2739_),
    .X(_2775_));
 sky130_fd_sc_hd__a2111o_1 _6154_ (.A1(\mem[25][8] ),
    .A2(_2736_),
    .B1(_2773_),
    .C1(_2774_),
    .D1(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__and3_1 _6155_ (.A(\mem[15][8] ),
    .B(_1435_),
    .C(_2592_),
    .X(_2777_));
 sky130_fd_sc_hd__and3_1 _6156_ (.A(\mem[24][8] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2778_));
 sky130_fd_sc_hd__and3_1 _6157_ (.A(\mem[13][8] ),
    .B(_1470_),
    .C(_2745_),
    .X(_2779_));
 sky130_fd_sc_hd__a2111o_1 _6158_ (.A1(\mem[10][8] ),
    .A2(_2742_),
    .B1(_2777_),
    .C1(_2778_),
    .D1(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__clkbuf_4 _6159_ (.A(_1034_),
    .X(_2781_));
 sky130_fd_sc_hd__inv_2 _6160_ (.A(\mem[19][8] ),
    .Y(_2782_));
 sky130_fd_sc_hd__or3_1 _6161_ (.A(_2782_),
    .B(_2598_),
    .C(_2655_),
    .X(_2783_));
 sky130_fd_sc_hd__or3b_1 _6162_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][8] ),
    .X(_2784_));
 sky130_fd_sc_hd__buf_2 _6163_ (.A(_1037_),
    .X(_2785_));
 sky130_fd_sc_hd__or3b_1 _6164_ (.A(_1445_),
    .B(_2785_),
    .C_N(\mem[1][8] ),
    .X(_2786_));
 sky130_fd_sc_hd__o2111ai_1 _6165_ (.A1(_1833_),
    .A2(_2781_),
    .B1(_2783_),
    .C1(_2784_),
    .D1(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__and3_1 _6166_ (.A(\mem[4][8] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2788_));
 sky130_fd_sc_hd__and3_1 _6167_ (.A(\mem[22][8] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2789_));
 sky130_fd_sc_hd__and3_1 _6168_ (.A(\mem[20][8] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2790_));
 sky130_fd_sc_hd__a2111o_1 _6169_ (.A1(\mem[18][8] ),
    .A2(_2753_),
    .B1(_2788_),
    .C1(_2789_),
    .D1(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__or4_1 _6170_ (.A(_2776_),
    .B(_2780_),
    .C(_2787_),
    .D(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__buf_4 _6171_ (.A(_1068_),
    .X(_2793_));
 sky130_fd_sc_hd__buf_4 _6172_ (.A(_1078_),
    .X(_2794_));
 sky130_fd_sc_hd__a22o_1 _6173_ (.A1(\mem[9][8] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][8] ),
    .X(_2795_));
 sky130_fd_sc_hd__buf_4 _6174_ (.A(_1070_),
    .X(_2796_));
 sky130_fd_sc_hd__a22o_1 _6175_ (.A1(\mem[27][8] ),
    .A2(_2796_),
    .B1(_1454_),
    .B2(\mem[28][8] ),
    .X(_2797_));
 sky130_fd_sc_hd__buf_4 _6176_ (.A(_1074_),
    .X(_2798_));
 sky130_fd_sc_hd__a32o_1 _6177_ (.A1(_2579_),
    .A2(\mem[31][8] ),
    .A3(_1456_),
    .B1(_2798_),
    .B2(\mem[14][8] ),
    .X(_2799_));
 sky130_fd_sc_hd__a2111o_1 _6178_ (.A1(\mem[26][8] ),
    .A2(_2793_),
    .B1(_2795_),
    .C1(_2797_),
    .D1(_2799_),
    .X(_2800_));
 sky130_fd_sc_hd__buf_4 _6179_ (.A(_1082_),
    .X(_2801_));
 sky130_fd_sc_hd__buf_4 _6180_ (.A(_1084_),
    .X(_2802_));
 sky130_fd_sc_hd__a22o_1 _6181_ (.A1(\mem[16][8] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][8] ),
    .X(_2803_));
 sky130_fd_sc_hd__a221o_1 _6182_ (.A1(\mem[8][8] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][8] ),
    .C1(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__clkbuf_8 _6183_ (.A(_1092_),
    .X(_2805_));
 sky130_fd_sc_hd__clkbuf_8 _6184_ (.A(_1094_),
    .X(_2806_));
 sky130_fd_sc_hd__buf_4 _6185_ (.A(_1096_),
    .X(_2807_));
 sky130_fd_sc_hd__clkbuf_8 _6186_ (.A(_1098_),
    .X(_2808_));
 sky130_fd_sc_hd__a22o_1 _6187_ (.A1(\mem[21][8] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][8] ),
    .X(_2809_));
 sky130_fd_sc_hd__a221o_1 _6188_ (.A1(\mem[2][8] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][8] ),
    .C1(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__or4_4 _6189_ (.A(_2792_),
    .B(_2800_),
    .C(_2804_),
    .D(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__clkbuf_1 _6190_ (.A(_2811_),
    .X(net112));
 sky130_fd_sc_hd__and3_1 _6191_ (.A(\mem[12][9] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2812_));
 sky130_fd_sc_hd__and3_1 _6192_ (.A(\mem[29][9] ),
    .B(_2588_),
    .C(_2705_),
    .X(_2813_));
 sky130_fd_sc_hd__and3_1 _6193_ (.A(\mem[30][9] ),
    .B(_2619_),
    .C(_2739_),
    .X(_2814_));
 sky130_fd_sc_hd__a2111o_1 _6194_ (.A1(\mem[25][9] ),
    .A2(_2736_),
    .B1(_2812_),
    .C1(_2813_),
    .D1(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__clkbuf_4 _6195_ (.A(_1018_),
    .X(_2816_));
 sky130_fd_sc_hd__and3_1 _6196_ (.A(\mem[15][9] ),
    .B(_2816_),
    .C(_2592_),
    .X(_2817_));
 sky130_fd_sc_hd__and3_1 _6197_ (.A(\mem[24][9] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2818_));
 sky130_fd_sc_hd__and3_1 _6198_ (.A(\mem[13][9] ),
    .B(_1470_),
    .C(_2745_),
    .X(_2819_));
 sky130_fd_sc_hd__a2111o_1 _6199_ (.A1(\mem[10][9] ),
    .A2(_2742_),
    .B1(_2817_),
    .C1(_2818_),
    .D1(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__inv_2 _6200_ (.A(\mem[19][9] ),
    .Y(_2821_));
 sky130_fd_sc_hd__or3_1 _6201_ (.A(_2821_),
    .B(_2598_),
    .C(_2655_),
    .X(_2822_));
 sky130_fd_sc_hd__or3b_1 _6202_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][9] ),
    .X(_2823_));
 sky130_fd_sc_hd__buf_2 _6203_ (.A(_1010_),
    .X(_2824_));
 sky130_fd_sc_hd__or3b_1 _6204_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][9] ),
    .X(_2825_));
 sky130_fd_sc_hd__o2111ai_1 _6205_ (.A1(_1864_),
    .A2(_2781_),
    .B1(_2822_),
    .C1(_2823_),
    .D1(_2825_),
    .Y(_2826_));
 sky130_fd_sc_hd__and3_1 _6206_ (.A(\mem[4][9] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2827_));
 sky130_fd_sc_hd__and3_1 _6207_ (.A(\mem[22][9] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2828_));
 sky130_fd_sc_hd__and3_1 _6208_ (.A(\mem[20][9] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2829_));
 sky130_fd_sc_hd__a2111o_1 _6209_ (.A1(\mem[18][9] ),
    .A2(_2753_),
    .B1(_2827_),
    .C1(_2828_),
    .D1(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__or4_1 _6210_ (.A(_2815_),
    .B(_2820_),
    .C(_2826_),
    .D(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__a22o_1 _6211_ (.A1(\mem[9][9] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][9] ),
    .X(_2832_));
 sky130_fd_sc_hd__buf_4 _6212_ (.A(_1071_),
    .X(_2833_));
 sky130_fd_sc_hd__a22o_1 _6213_ (.A1(\mem[27][9] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][9] ),
    .X(_2834_));
 sky130_fd_sc_hd__buf_4 _6214_ (.A(_1028_),
    .X(_2835_));
 sky130_fd_sc_hd__a32o_1 _6215_ (.A1(_2579_),
    .A2(\mem[31][9] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][9] ),
    .X(_2836_));
 sky130_fd_sc_hd__a2111o_1 _6216_ (.A1(\mem[26][9] ),
    .A2(_2793_),
    .B1(_2832_),
    .C1(_2834_),
    .D1(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__a22o_1 _6217_ (.A1(\mem[16][9] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][9] ),
    .X(_2838_));
 sky130_fd_sc_hd__a221o_1 _6218_ (.A1(\mem[8][9] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][9] ),
    .C1(_2838_),
    .X(_2839_));
 sky130_fd_sc_hd__a22o_1 _6219_ (.A1(\mem[21][9] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][9] ),
    .X(_2840_));
 sky130_fd_sc_hd__a221o_1 _6220_ (.A1(\mem[2][9] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][9] ),
    .C1(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__or4_4 _6221_ (.A(_2831_),
    .B(_2837_),
    .C(_2839_),
    .D(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__clkbuf_1 _6222_ (.A(_2842_),
    .X(net113));
 sky130_fd_sc_hd__and3_1 _6223_ (.A(\mem[12][10] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2843_));
 sky130_fd_sc_hd__and3_1 _6224_ (.A(\mem[29][10] ),
    .B(_2588_),
    .C(_2705_),
    .X(_2844_));
 sky130_fd_sc_hd__and3_1 _6225_ (.A(\mem[30][10] ),
    .B(_2619_),
    .C(_2739_),
    .X(_2845_));
 sky130_fd_sc_hd__a2111o_1 _6226_ (.A1(\mem[25][10] ),
    .A2(_2736_),
    .B1(_2843_),
    .C1(_2844_),
    .D1(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__and3_1 _6227_ (.A(\mem[15][10] ),
    .B(_2816_),
    .C(_2592_),
    .X(_2847_));
 sky130_fd_sc_hd__and3_1 _6228_ (.A(\mem[24][10] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2848_));
 sky130_fd_sc_hd__and3_1 _6229_ (.A(\mem[13][10] ),
    .B(_1019_),
    .C(_2745_),
    .X(_2849_));
 sky130_fd_sc_hd__a2111o_1 _6230_ (.A1(\mem[10][10] ),
    .A2(_2742_),
    .B1(_2847_),
    .C1(_2848_),
    .D1(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__clkinv_2 _6231_ (.A(\mem[19][10] ),
    .Y(_2851_));
 sky130_fd_sc_hd__or3_1 _6232_ (.A(_2851_),
    .B(_2598_),
    .C(_2655_),
    .X(_2852_));
 sky130_fd_sc_hd__or3b_1 _6233_ (.A(_2568_),
    .B(_1443_),
    .C_N(\mem[5][10] ),
    .X(_2853_));
 sky130_fd_sc_hd__or3b_1 _6234_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][10] ),
    .X(_2854_));
 sky130_fd_sc_hd__o2111ai_1 _6235_ (.A1(_1896_),
    .A2(_2781_),
    .B1(_2852_),
    .C1(_2853_),
    .D1(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__and3_1 _6236_ (.A(\mem[4][10] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2856_));
 sky130_fd_sc_hd__and3_1 _6237_ (.A(\mem[22][10] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2857_));
 sky130_fd_sc_hd__and3_1 _6238_ (.A(\mem[20][10] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2858_));
 sky130_fd_sc_hd__a2111o_1 _6239_ (.A1(\mem[18][10] ),
    .A2(_2753_),
    .B1(_2856_),
    .C1(_2857_),
    .D1(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__or4_1 _6240_ (.A(_2846_),
    .B(_2850_),
    .C(_2855_),
    .D(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__a22o_1 _6241_ (.A1(\mem[9][10] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][10] ),
    .X(_2861_));
 sky130_fd_sc_hd__a22o_1 _6242_ (.A1(\mem[27][10] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][10] ),
    .X(_2862_));
 sky130_fd_sc_hd__a32o_1 _6243_ (.A1(_2579_),
    .A2(\mem[31][10] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][10] ),
    .X(_2863_));
 sky130_fd_sc_hd__a2111o_1 _6244_ (.A1(\mem[26][10] ),
    .A2(_2793_),
    .B1(_2861_),
    .C1(_2862_),
    .D1(_2863_),
    .X(_2864_));
 sky130_fd_sc_hd__a22o_1 _6245_ (.A1(\mem[16][10] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][10] ),
    .X(_2865_));
 sky130_fd_sc_hd__a221o_1 _6246_ (.A1(\mem[8][10] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][10] ),
    .C1(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__a22o_1 _6247_ (.A1(\mem[21][10] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][10] ),
    .X(_2867_));
 sky130_fd_sc_hd__a221o_1 _6248_ (.A1(\mem[2][10] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][10] ),
    .C1(_2867_),
    .X(_2868_));
 sky130_fd_sc_hd__or4_1 _6249_ (.A(_2860_),
    .B(_2864_),
    .C(_2866_),
    .D(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__buf_8 _6250_ (.A(_2869_),
    .X(net83));
 sky130_fd_sc_hd__and3_1 _6251_ (.A(\mem[12][11] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2870_));
 sky130_fd_sc_hd__and3_1 _6252_ (.A(\mem[29][11] ),
    .B(_2588_),
    .C(_2705_),
    .X(_2871_));
 sky130_fd_sc_hd__and3_1 _6253_ (.A(\mem[30][11] ),
    .B(_2619_),
    .C(_2739_),
    .X(_2872_));
 sky130_fd_sc_hd__a2111o_1 _6254_ (.A1(\mem[25][11] ),
    .A2(_2736_),
    .B1(_2870_),
    .C1(_2871_),
    .D1(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__and3_1 _6255_ (.A(\mem[15][11] ),
    .B(_2816_),
    .C(_2592_),
    .X(_2874_));
 sky130_fd_sc_hd__and3_1 _6256_ (.A(\mem[24][11] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2875_));
 sky130_fd_sc_hd__and3_1 _6257_ (.A(\mem[13][11] ),
    .B(_1019_),
    .C(_2745_),
    .X(_2876_));
 sky130_fd_sc_hd__a2111o_1 _6258_ (.A1(\mem[10][11] ),
    .A2(_2742_),
    .B1(_2874_),
    .C1(_2875_),
    .D1(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__inv_2 _6259_ (.A(\mem[19][11] ),
    .Y(_2878_));
 sky130_fd_sc_hd__or3_1 _6260_ (.A(_2878_),
    .B(_2598_),
    .C(_2655_),
    .X(_2879_));
 sky130_fd_sc_hd__or3b_1 _6261_ (.A(_2568_),
    .B(_1180_),
    .C_N(\mem[5][11] ),
    .X(_2880_));
 sky130_fd_sc_hd__or3b_1 _6262_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][11] ),
    .X(_2881_));
 sky130_fd_sc_hd__o2111ai_1 _6263_ (.A1(_1934_),
    .A2(_2781_),
    .B1(_2879_),
    .C1(_2880_),
    .D1(_2881_),
    .Y(_2882_));
 sky130_fd_sc_hd__and3_1 _6264_ (.A(\mem[4][11] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2883_));
 sky130_fd_sc_hd__and3_1 _6265_ (.A(\mem[22][11] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2884_));
 sky130_fd_sc_hd__and3_1 _6266_ (.A(\mem[20][11] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2885_));
 sky130_fd_sc_hd__a2111o_1 _6267_ (.A1(\mem[18][11] ),
    .A2(_2753_),
    .B1(_2883_),
    .C1(_2884_),
    .D1(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__or4_1 _6268_ (.A(_2873_),
    .B(_2877_),
    .C(_2882_),
    .D(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__a22o_1 _6269_ (.A1(\mem[9][11] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][11] ),
    .X(_2888_));
 sky130_fd_sc_hd__a22o_1 _6270_ (.A1(\mem[27][11] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][11] ),
    .X(_2889_));
 sky130_fd_sc_hd__a32o_1 _6271_ (.A1(_1131_),
    .A2(\mem[31][11] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][11] ),
    .X(_2890_));
 sky130_fd_sc_hd__a2111o_1 _6272_ (.A1(\mem[26][11] ),
    .A2(_2793_),
    .B1(_2888_),
    .C1(_2889_),
    .D1(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__a22o_1 _6273_ (.A1(\mem[16][11] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][11] ),
    .X(_2892_));
 sky130_fd_sc_hd__a221o_1 _6274_ (.A1(\mem[8][11] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][11] ),
    .C1(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__a22o_1 _6275_ (.A1(\mem[21][11] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][11] ),
    .X(_2894_));
 sky130_fd_sc_hd__a221o_1 _6276_ (.A1(\mem[2][11] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][11] ),
    .C1(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__or4_4 _6277_ (.A(_2887_),
    .B(_2891_),
    .C(_2893_),
    .D(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__clkbuf_1 _6278_ (.A(_2896_),
    .X(net84));
 sky130_fd_sc_hd__and3_1 _6279_ (.A(\mem[12][12] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2897_));
 sky130_fd_sc_hd__and3_1 _6280_ (.A(\mem[29][12] ),
    .B(_1067_),
    .C(_2705_),
    .X(_2898_));
 sky130_fd_sc_hd__and3_1 _6281_ (.A(\mem[30][12] ),
    .B(_2619_),
    .C(_2739_),
    .X(_2899_));
 sky130_fd_sc_hd__a2111o_1 _6282_ (.A1(\mem[25][12] ),
    .A2(_2736_),
    .B1(_2897_),
    .C1(_2898_),
    .D1(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__and3_1 _6283_ (.A(\mem[15][12] ),
    .B(_2816_),
    .C(_1027_),
    .X(_2901_));
 sky130_fd_sc_hd__and3_1 _6284_ (.A(\mem[24][12] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2902_));
 sky130_fd_sc_hd__and3_1 _6285_ (.A(\mem[13][12] ),
    .B(_1019_),
    .C(_2745_),
    .X(_2903_));
 sky130_fd_sc_hd__a2111o_1 _6286_ (.A1(\mem[10][12] ),
    .A2(_2742_),
    .B1(_2901_),
    .C1(_2902_),
    .D1(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__or3b_1 _6287_ (.A(_1057_),
    .B(_1040_),
    .C_N(\mem[5][12] ),
    .X(_2905_));
 sky130_fd_sc_hd__inv_2 _6288_ (.A(\mem[19][12] ),
    .Y(_2906_));
 sky130_fd_sc_hd__or3_1 _6289_ (.A(_2906_),
    .B(_1045_),
    .C(_1046_),
    .X(_2907_));
 sky130_fd_sc_hd__or3b_1 _6290_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][12] ),
    .X(_2908_));
 sky130_fd_sc_hd__o2111ai_1 _6291_ (.A1(_1971_),
    .A2(_2781_),
    .B1(_2905_),
    .C1(_2907_),
    .D1(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__and3_1 _6292_ (.A(\mem[4][12] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2910_));
 sky130_fd_sc_hd__and3_1 _6293_ (.A(\mem[22][12] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2911_));
 sky130_fd_sc_hd__and3_1 _6294_ (.A(\mem[20][12] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2912_));
 sky130_fd_sc_hd__a2111o_1 _6295_ (.A1(\mem[18][12] ),
    .A2(_2753_),
    .B1(_2910_),
    .C1(_2911_),
    .D1(_2912_),
    .X(_2913_));
 sky130_fd_sc_hd__or4_1 _6296_ (.A(_2900_),
    .B(_2904_),
    .C(_2909_),
    .D(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__a22o_1 _6297_ (.A1(\mem[9][12] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][12] ),
    .X(_2915_));
 sky130_fd_sc_hd__a22o_1 _6298_ (.A1(\mem[27][12] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][12] ),
    .X(_2916_));
 sky130_fd_sc_hd__a32o_1 _6299_ (.A1(_1131_),
    .A2(\mem[31][12] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][12] ),
    .X(_2917_));
 sky130_fd_sc_hd__a2111o_1 _6300_ (.A1(\mem[26][12] ),
    .A2(_2793_),
    .B1(_2915_),
    .C1(_2916_),
    .D1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__a22o_1 _6301_ (.A1(\mem[16][12] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][12] ),
    .X(_2919_));
 sky130_fd_sc_hd__a221o_1 _6302_ (.A1(\mem[8][12] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][12] ),
    .C1(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__a22o_1 _6303_ (.A1(\mem[21][12] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][12] ),
    .X(_2921_));
 sky130_fd_sc_hd__a221o_1 _6304_ (.A1(\mem[2][12] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][12] ),
    .C1(_2921_),
    .X(_2922_));
 sky130_fd_sc_hd__or4_1 _6305_ (.A(_2914_),
    .B(_2918_),
    .C(_2920_),
    .D(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__clkbuf_4 _6306_ (.A(_2923_),
    .X(net85));
 sky130_fd_sc_hd__and3_1 _6307_ (.A(\mem[12][13] ),
    .B(_2703_),
    .C(_2645_),
    .X(_2924_));
 sky130_fd_sc_hd__and3_1 _6308_ (.A(\mem[29][13] ),
    .B(_1067_),
    .C(_2705_),
    .X(_2925_));
 sky130_fd_sc_hd__and3_1 _6309_ (.A(\mem[30][13] ),
    .B(_1006_),
    .C(_2739_),
    .X(_2926_));
 sky130_fd_sc_hd__a2111o_1 _6310_ (.A1(\mem[25][13] ),
    .A2(_2736_),
    .B1(_2924_),
    .C1(_2925_),
    .D1(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__and3_1 _6311_ (.A(\mem[15][13] ),
    .B(_2816_),
    .C(_1027_),
    .X(_2928_));
 sky130_fd_sc_hd__and3_1 _6312_ (.A(\mem[24][13] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2929_));
 sky130_fd_sc_hd__and3_1 _6313_ (.A(\mem[13][13] ),
    .B(_1019_),
    .C(_2745_),
    .X(_2930_));
 sky130_fd_sc_hd__a2111o_1 _6314_ (.A1(\mem[10][13] ),
    .A2(_2742_),
    .B1(_2928_),
    .C1(_2929_),
    .D1(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__inv_2 _6315_ (.A(\mem[19][13] ),
    .Y(_2932_));
 sky130_fd_sc_hd__or3_1 _6316_ (.A(_2932_),
    .B(_2598_),
    .C(_2655_),
    .X(_2933_));
 sky130_fd_sc_hd__or3b_1 _6317_ (.A(_2568_),
    .B(_1180_),
    .C_N(\mem[5][13] ),
    .X(_2934_));
 sky130_fd_sc_hd__or3b_1 _6318_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][13] ),
    .X(_2935_));
 sky130_fd_sc_hd__o2111ai_1 _6319_ (.A1(_1998_),
    .A2(_2781_),
    .B1(_2933_),
    .C1(_2934_),
    .D1(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__and3_1 _6320_ (.A(\mem[4][13] ),
    .B(_2719_),
    .C(_2660_),
    .X(_2937_));
 sky130_fd_sc_hd__and3_1 _6321_ (.A(\mem[22][13] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2938_));
 sky130_fd_sc_hd__and3_1 _6322_ (.A(\mem[20][13] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2939_));
 sky130_fd_sc_hd__a2111o_1 _6323_ (.A1(\mem[18][13] ),
    .A2(_2753_),
    .B1(_2937_),
    .C1(_2938_),
    .D1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__or4_1 _6324_ (.A(_2927_),
    .B(_2931_),
    .C(_2936_),
    .D(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__a22o_1 _6325_ (.A1(\mem[9][13] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][13] ),
    .X(_2942_));
 sky130_fd_sc_hd__a22o_1 _6326_ (.A1(\mem[27][13] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][13] ),
    .X(_2943_));
 sky130_fd_sc_hd__a32o_1 _6327_ (.A1(_1131_),
    .A2(\mem[31][13] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][13] ),
    .X(_2944_));
 sky130_fd_sc_hd__a2111o_1 _6328_ (.A1(\mem[26][13] ),
    .A2(_2793_),
    .B1(_2942_),
    .C1(_2943_),
    .D1(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__a22o_1 _6329_ (.A1(\mem[16][13] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][13] ),
    .X(_2946_));
 sky130_fd_sc_hd__a221o_1 _6330_ (.A1(\mem[8][13] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][13] ),
    .C1(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__a22o_1 _6331_ (.A1(\mem[21][13] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][13] ),
    .X(_2948_));
 sky130_fd_sc_hd__a221o_1 _6332_ (.A1(\mem[2][13] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][13] ),
    .C1(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__or4_1 _6333_ (.A(_2941_),
    .B(_2945_),
    .C(_2947_),
    .D(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__clkbuf_2 _6334_ (.A(_2950_),
    .X(net86));
 sky130_fd_sc_hd__and3_1 _6335_ (.A(\mem[12][14] ),
    .B(_2703_),
    .C(_1003_),
    .X(_2951_));
 sky130_fd_sc_hd__and3_1 _6336_ (.A(\mem[29][14] ),
    .B(_1067_),
    .C(_2705_),
    .X(_2952_));
 sky130_fd_sc_hd__and3_1 _6337_ (.A(\mem[30][14] ),
    .B(_1006_),
    .C(_2739_),
    .X(_2953_));
 sky130_fd_sc_hd__a2111o_1 _6338_ (.A1(\mem[25][14] ),
    .A2(_2736_),
    .B1(_2951_),
    .C1(_2952_),
    .D1(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__and3_1 _6339_ (.A(\mem[15][14] ),
    .B(_2816_),
    .C(_1027_),
    .X(_2955_));
 sky130_fd_sc_hd__and3_1 _6340_ (.A(\mem[24][14] ),
    .B(_2710_),
    .C(_2680_),
    .X(_2956_));
 sky130_fd_sc_hd__and3_1 _6341_ (.A(\mem[13][14] ),
    .B(_1019_),
    .C(_2745_),
    .X(_2957_));
 sky130_fd_sc_hd__a2111o_1 _6342_ (.A1(\mem[10][14] ),
    .A2(_2742_),
    .B1(_2955_),
    .C1(_2956_),
    .D1(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__inv_2 _6343_ (.A(\mem[19][14] ),
    .Y(_2959_));
 sky130_fd_sc_hd__or3_1 _6344_ (.A(_2959_),
    .B(_2598_),
    .C(_2655_),
    .X(_2960_));
 sky130_fd_sc_hd__or3b_1 _6345_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][14] ),
    .X(_2961_));
 sky130_fd_sc_hd__or3b_1 _6346_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][14] ),
    .X(_2962_));
 sky130_fd_sc_hd__o2111ai_1 _6347_ (.A1(_2025_),
    .A2(_2781_),
    .B1(_2960_),
    .C1(_2961_),
    .D1(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__and3_1 _6348_ (.A(\mem[4][14] ),
    .B(_2719_),
    .C(_1054_),
    .X(_2964_));
 sky130_fd_sc_hd__and3_1 _6349_ (.A(\mem[22][14] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2965_));
 sky130_fd_sc_hd__and3_1 _6350_ (.A(\mem[20][14] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2966_));
 sky130_fd_sc_hd__a2111o_1 _6351_ (.A1(\mem[18][14] ),
    .A2(_2753_),
    .B1(_2964_),
    .C1(_2965_),
    .D1(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__or4_1 _6352_ (.A(_2954_),
    .B(_2958_),
    .C(_2963_),
    .D(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__a22o_1 _6353_ (.A1(\mem[9][14] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][14] ),
    .X(_2969_));
 sky130_fd_sc_hd__a22o_1 _6354_ (.A1(\mem[27][14] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][14] ),
    .X(_2970_));
 sky130_fd_sc_hd__a32o_1 _6355_ (.A1(_1131_),
    .A2(\mem[31][14] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][14] ),
    .X(_2971_));
 sky130_fd_sc_hd__a2111o_1 _6356_ (.A1(\mem[26][14] ),
    .A2(_2793_),
    .B1(_2969_),
    .C1(_2970_),
    .D1(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__a22o_1 _6357_ (.A1(\mem[16][14] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][14] ),
    .X(_2973_));
 sky130_fd_sc_hd__a221o_1 _6358_ (.A1(\mem[8][14] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][14] ),
    .C1(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__a22o_1 _6359_ (.A1(\mem[21][14] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][14] ),
    .X(_2975_));
 sky130_fd_sc_hd__a221o_1 _6360_ (.A1(\mem[2][14] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][14] ),
    .C1(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__or4_4 _6361_ (.A(_2968_),
    .B(_2972_),
    .C(_2974_),
    .D(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__clkbuf_1 _6362_ (.A(_2977_),
    .X(net87));
 sky130_fd_sc_hd__and3_1 _6363_ (.A(\mem[12][15] ),
    .B(_2703_),
    .C(_1003_),
    .X(_2978_));
 sky130_fd_sc_hd__and3_1 _6364_ (.A(\mem[29][15] ),
    .B(_1067_),
    .C(_2705_),
    .X(_2979_));
 sky130_fd_sc_hd__and3_1 _6365_ (.A(\mem[30][15] ),
    .B(_1006_),
    .C(_2739_),
    .X(_2980_));
 sky130_fd_sc_hd__a2111o_1 _6366_ (.A1(\mem[25][15] ),
    .A2(_2736_),
    .B1(_2978_),
    .C1(_2979_),
    .D1(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__and3_1 _6367_ (.A(\mem[15][15] ),
    .B(_2816_),
    .C(_1027_),
    .X(_2982_));
 sky130_fd_sc_hd__and3_1 _6368_ (.A(\mem[24][15] ),
    .B(_2710_),
    .C(_1062_),
    .X(_2983_));
 sky130_fd_sc_hd__and3_1 _6369_ (.A(\mem[13][15] ),
    .B(_1019_),
    .C(_2745_),
    .X(_2984_));
 sky130_fd_sc_hd__a2111o_1 _6370_ (.A1(\mem[10][15] ),
    .A2(_2742_),
    .B1(_2982_),
    .C1(_2983_),
    .D1(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__inv_2 _6371_ (.A(\mem[19][15] ),
    .Y(_2986_));
 sky130_fd_sc_hd__or3_1 _6372_ (.A(_2986_),
    .B(_1026_),
    .C(_2655_),
    .X(_2987_));
 sky130_fd_sc_hd__or3b_1 _6373_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][15] ),
    .X(_2988_));
 sky130_fd_sc_hd__or3b_1 _6374_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][15] ),
    .X(_2989_));
 sky130_fd_sc_hd__o2111ai_1 _6375_ (.A1(_2056_),
    .A2(_2781_),
    .B1(_2987_),
    .C1(_2988_),
    .D1(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__and3_1 _6376_ (.A(\mem[4][15] ),
    .B(_2719_),
    .C(_1054_),
    .X(_2991_));
 sky130_fd_sc_hd__and3_1 _6377_ (.A(\mem[22][15] ),
    .B(_2721_),
    .C(_2722_),
    .X(_2992_));
 sky130_fd_sc_hd__and3_1 _6378_ (.A(\mem[20][15] ),
    .B(_2756_),
    .C(_2757_),
    .X(_2993_));
 sky130_fd_sc_hd__a2111o_1 _6379_ (.A1(\mem[18][15] ),
    .A2(_2753_),
    .B1(_2991_),
    .C1(_2992_),
    .D1(_2993_),
    .X(_2994_));
 sky130_fd_sc_hd__or4_1 _6380_ (.A(_2981_),
    .B(_2985_),
    .C(_2990_),
    .D(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__a22o_1 _6381_ (.A1(\mem[9][15] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][15] ),
    .X(_2996_));
 sky130_fd_sc_hd__a22o_1 _6382_ (.A1(\mem[27][15] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][15] ),
    .X(_2997_));
 sky130_fd_sc_hd__a32o_1 _6383_ (.A1(_1131_),
    .A2(\mem[31][15] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][15] ),
    .X(_2998_));
 sky130_fd_sc_hd__a2111o_1 _6384_ (.A1(\mem[26][15] ),
    .A2(_2793_),
    .B1(_2996_),
    .C1(_2997_),
    .D1(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__a22o_1 _6385_ (.A1(\mem[16][15] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][15] ),
    .X(_3000_));
 sky130_fd_sc_hd__a221o_1 _6386_ (.A1(\mem[8][15] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][15] ),
    .C1(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__a22o_1 _6387_ (.A1(\mem[21][15] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][15] ),
    .X(_3002_));
 sky130_fd_sc_hd__a221o_1 _6388_ (.A1(\mem[2][15] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][15] ),
    .C1(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__or4_1 _6389_ (.A(_2995_),
    .B(_2999_),
    .C(_3001_),
    .D(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__buf_2 _6390_ (.A(_3004_),
    .X(net88));
 sky130_fd_sc_hd__and3_1 _6391_ (.A(\mem[12][16] ),
    .B(_1000_),
    .C(_1003_),
    .X(_3005_));
 sky130_fd_sc_hd__and3_1 _6392_ (.A(\mem[29][16] ),
    .B(_1067_),
    .C(_1007_),
    .X(_3006_));
 sky130_fd_sc_hd__and3_1 _6393_ (.A(\mem[30][16] ),
    .B(_1006_),
    .C(_2739_),
    .X(_3007_));
 sky130_fd_sc_hd__a2111o_1 _6394_ (.A1(\mem[25][16] ),
    .A2(_2736_),
    .B1(_3005_),
    .C1(_3006_),
    .D1(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__and3_1 _6395_ (.A(\mem[15][16] ),
    .B(_2816_),
    .C(_1027_),
    .X(_3009_));
 sky130_fd_sc_hd__and3_1 _6396_ (.A(\mem[24][16] ),
    .B(_1021_),
    .C(_1062_),
    .X(_3010_));
 sky130_fd_sc_hd__and3_1 _6397_ (.A(\mem[13][16] ),
    .B(_1019_),
    .C(_2745_),
    .X(_3011_));
 sky130_fd_sc_hd__a2111o_1 _6398_ (.A1(\mem[10][16] ),
    .A2(_2742_),
    .B1(_3009_),
    .C1(_3010_),
    .D1(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__inv_2 _6399_ (.A(\mem[19][16] ),
    .Y(_3013_));
 sky130_fd_sc_hd__or3_1 _6400_ (.A(_3013_),
    .B(_1026_),
    .C(_1032_),
    .X(_3014_));
 sky130_fd_sc_hd__or3b_1 _6401_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][16] ),
    .X(_3015_));
 sky130_fd_sc_hd__or3b_1 _6402_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][16] ),
    .X(_3016_));
 sky130_fd_sc_hd__o2111ai_1 _6403_ (.A1(_2082_),
    .A2(_2781_),
    .B1(_3014_),
    .C1(_3015_),
    .D1(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__and3_1 _6404_ (.A(\mem[4][16] ),
    .B(_1004_),
    .C(_1054_),
    .X(_3018_));
 sky130_fd_sc_hd__and3_1 _6405_ (.A(\mem[22][16] ),
    .B(_1011_),
    .C(_1058_),
    .X(_3019_));
 sky130_fd_sc_hd__and3_1 _6406_ (.A(\mem[20][16] ),
    .B(_2756_),
    .C(_2757_),
    .X(_3020_));
 sky130_fd_sc_hd__a2111o_1 _6407_ (.A1(\mem[18][16] ),
    .A2(_2753_),
    .B1(_3018_),
    .C1(_3019_),
    .D1(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__or4_1 _6408_ (.A(_3008_),
    .B(_3012_),
    .C(_3017_),
    .D(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__a22o_1 _6409_ (.A1(\mem[9][16] ),
    .A2(_2761_),
    .B1(_2794_),
    .B2(\mem[11][16] ),
    .X(_3023_));
 sky130_fd_sc_hd__a22o_1 _6410_ (.A1(\mem[27][16] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][16] ),
    .X(_3024_));
 sky130_fd_sc_hd__a32o_1 _6411_ (.A1(_1131_),
    .A2(\mem[31][16] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][16] ),
    .X(_3025_));
 sky130_fd_sc_hd__a2111o_1 _6412_ (.A1(\mem[26][16] ),
    .A2(_2793_),
    .B1(_3023_),
    .C1(_3024_),
    .D1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__a22o_1 _6413_ (.A1(\mem[16][16] ),
    .A2(_2766_),
    .B1(_2767_),
    .B2(\mem[7][16] ),
    .X(_3027_));
 sky130_fd_sc_hd__a221o_1 _6414_ (.A1(\mem[8][16] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][16] ),
    .C1(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__a22o_1 _6415_ (.A1(\mem[21][16] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][16] ),
    .X(_3029_));
 sky130_fd_sc_hd__a221o_1 _6416_ (.A1(\mem[2][16] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][16] ),
    .C1(_3029_),
    .X(_3030_));
 sky130_fd_sc_hd__or4_2 _6417_ (.A(_3022_),
    .B(_3026_),
    .C(_3028_),
    .D(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__clkbuf_2 _6418_ (.A(_3031_),
    .X(net89));
 sky130_fd_sc_hd__and3_1 _6419_ (.A(\mem[12][17] ),
    .B(_1000_),
    .C(_1003_),
    .X(_3032_));
 sky130_fd_sc_hd__and3_1 _6420_ (.A(\mem[29][17] ),
    .B(_1067_),
    .C(_1007_),
    .X(_3033_));
 sky130_fd_sc_hd__and3_1 _6421_ (.A(\mem[30][17] ),
    .B(_1006_),
    .C(_1012_),
    .X(_3034_));
 sky130_fd_sc_hd__a2111o_1 _6422_ (.A1(\mem[25][17] ),
    .A2(_0996_),
    .B1(_3032_),
    .C1(_3033_),
    .D1(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__and3_1 _6423_ (.A(\mem[15][17] ),
    .B(_2816_),
    .C(_1027_),
    .X(_3036_));
 sky130_fd_sc_hd__and3_1 _6424_ (.A(\mem[24][17] ),
    .B(_1021_),
    .C(_1062_),
    .X(_3037_));
 sky130_fd_sc_hd__and3_1 _6425_ (.A(\mem[13][17] ),
    .B(_1019_),
    .C(_1008_),
    .X(_3038_));
 sky130_fd_sc_hd__a2111o_1 _6426_ (.A1(\mem[10][17] ),
    .A2(_1016_),
    .B1(_3036_),
    .C1(_3037_),
    .D1(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__inv_2 _6427_ (.A(\mem[19][17] ),
    .Y(_3040_));
 sky130_fd_sc_hd__or3_1 _6428_ (.A(_3040_),
    .B(_1026_),
    .C(_1032_),
    .X(_3041_));
 sky130_fd_sc_hd__or3b_1 _6429_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][17] ),
    .X(_3042_));
 sky130_fd_sc_hd__or3b_1 _6430_ (.A(_2824_),
    .B(_2785_),
    .C_N(\mem[1][17] ),
    .X(_3043_));
 sky130_fd_sc_hd__o2111ai_1 _6431_ (.A1(_2110_),
    .A2(_2781_),
    .B1(_3041_),
    .C1(_3042_),
    .D1(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__and3_1 _6432_ (.A(\mem[4][17] ),
    .B(_1004_),
    .C(_1054_),
    .X(_3045_));
 sky130_fd_sc_hd__and3_1 _6433_ (.A(\mem[22][17] ),
    .B(_1011_),
    .C(_1058_),
    .X(_3046_));
 sky130_fd_sc_hd__and3_1 _6434_ (.A(\mem[20][17] ),
    .B(_1055_),
    .C(_1024_),
    .X(_3047_));
 sky130_fd_sc_hd__a2111o_1 _6435_ (.A1(\mem[18][17] ),
    .A2(_1050_),
    .B1(_3045_),
    .C1(_3046_),
    .D1(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__or4_1 _6436_ (.A(_3035_),
    .B(_3039_),
    .C(_3044_),
    .D(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__a22o_1 _6437_ (.A1(\mem[9][17] ),
    .A2(_1076_),
    .B1(_2794_),
    .B2(\mem[11][17] ),
    .X(_3050_));
 sky130_fd_sc_hd__a22o_1 _6438_ (.A1(\mem[27][17] ),
    .A2(_2796_),
    .B1(_2833_),
    .B2(\mem[28][17] ),
    .X(_3051_));
 sky130_fd_sc_hd__a32o_1 _6439_ (.A1(_1131_),
    .A2(\mem[31][17] ),
    .A3(_2835_),
    .B1(_2798_),
    .B2(\mem[14][17] ),
    .X(_3052_));
 sky130_fd_sc_hd__a2111o_1 _6440_ (.A1(\mem[26][17] ),
    .A2(_2793_),
    .B1(_3050_),
    .C1(_3051_),
    .D1(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__a22o_1 _6441_ (.A1(\mem[16][17] ),
    .A2(_1086_),
    .B1(_1088_),
    .B2(\mem[7][17] ),
    .X(_3054_));
 sky130_fd_sc_hd__a221o_1 _6442_ (.A1(\mem[8][17] ),
    .A2(_2801_),
    .B1(_2802_),
    .B2(\mem[6][17] ),
    .C1(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__a22o_1 _6443_ (.A1(\mem[21][17] ),
    .A2(_2807_),
    .B1(_2808_),
    .B2(\mem[17][17] ),
    .X(_3056_));
 sky130_fd_sc_hd__a221o_1 _6444_ (.A1(\mem[2][17] ),
    .A2(_2805_),
    .B1(_2806_),
    .B2(\mem[23][17] ),
    .C1(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__or4_4 _6445_ (.A(_3049_),
    .B(_3053_),
    .C(_3055_),
    .D(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__clkbuf_1 _6446_ (.A(_3058_),
    .X(net90));
 sky130_fd_sc_hd__and3_1 _6447_ (.A(\mem[12][18] ),
    .B(_1000_),
    .C(_1003_),
    .X(_3059_));
 sky130_fd_sc_hd__and3_1 _6448_ (.A(\mem[29][18] ),
    .B(_1067_),
    .C(_1007_),
    .X(_3060_));
 sky130_fd_sc_hd__and3_1 _6449_ (.A(\mem[30][18] ),
    .B(_1006_),
    .C(_1012_),
    .X(_3061_));
 sky130_fd_sc_hd__a2111o_1 _6450_ (.A1(\mem[25][18] ),
    .A2(_0996_),
    .B1(_3059_),
    .C1(_3060_),
    .D1(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__and3_1 _6451_ (.A(\mem[15][18] ),
    .B(_2816_),
    .C(_1027_),
    .X(_3063_));
 sky130_fd_sc_hd__and3_1 _6452_ (.A(\mem[24][18] ),
    .B(_1021_),
    .C(_1062_),
    .X(_3064_));
 sky130_fd_sc_hd__and3_1 _6453_ (.A(\mem[13][18] ),
    .B(_1019_),
    .C(_1008_),
    .X(_3065_));
 sky130_fd_sc_hd__a2111o_1 _6454_ (.A1(\mem[10][18] ),
    .A2(_1016_),
    .B1(_3063_),
    .C1(_3064_),
    .D1(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__clkinv_2 _6455_ (.A(\mem[19][18] ),
    .Y(_3067_));
 sky130_fd_sc_hd__or3_1 _6456_ (.A(_3067_),
    .B(_1026_),
    .C(_1032_),
    .X(_3068_));
 sky130_fd_sc_hd__or3b_1 _6457_ (.A(_1036_),
    .B(_1180_),
    .C_N(\mem[5][18] ),
    .X(_3069_));
 sky130_fd_sc_hd__or3b_1 _6458_ (.A(_2824_),
    .B(_1037_),
    .C_N(\mem[1][18] ),
    .X(_3070_));
 sky130_fd_sc_hd__o2111ai_1 _6459_ (.A1(_2141_),
    .A2(_1034_),
    .B1(_3068_),
    .C1(_3069_),
    .D1(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__and3_1 _6460_ (.A(\mem[4][18] ),
    .B(_1004_),
    .C(_1054_),
    .X(_3072_));
 sky130_fd_sc_hd__and3_1 _6461_ (.A(\mem[22][18] ),
    .B(_1011_),
    .C(_1058_),
    .X(_3073_));
 sky130_fd_sc_hd__and3_1 _6462_ (.A(\mem[20][18] ),
    .B(_1055_),
    .C(_1024_),
    .X(_3074_));
 sky130_fd_sc_hd__a2111o_1 _6463_ (.A1(\mem[18][18] ),
    .A2(_1050_),
    .B1(_3072_),
    .C1(_3073_),
    .D1(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__or4_1 _6464_ (.A(_3062_),
    .B(_3066_),
    .C(_3071_),
    .D(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__a22o_1 _6465_ (.A1(\mem[9][18] ),
    .A2(_1076_),
    .B1(_1078_),
    .B2(\mem[11][18] ),
    .X(_3077_));
 sky130_fd_sc_hd__a22o_1 _6466_ (.A1(\mem[27][18] ),
    .A2(_1070_),
    .B1(_2833_),
    .B2(\mem[28][18] ),
    .X(_3078_));
 sky130_fd_sc_hd__a32o_1 _6467_ (.A1(_1131_),
    .A2(\mem[31][18] ),
    .A3(_2835_),
    .B1(_1074_),
    .B2(\mem[14][18] ),
    .X(_3079_));
 sky130_fd_sc_hd__a2111o_1 _6468_ (.A1(\mem[26][18] ),
    .A2(_1068_),
    .B1(_3077_),
    .C1(_3078_),
    .D1(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__a22o_1 _6469_ (.A1(\mem[16][18] ),
    .A2(_1086_),
    .B1(_1088_),
    .B2(\mem[7][18] ),
    .X(_3081_));
 sky130_fd_sc_hd__a221o_1 _6470_ (.A1(\mem[8][18] ),
    .A2(_1082_),
    .B1(_1084_),
    .B2(\mem[6][18] ),
    .C1(_3081_),
    .X(_3082_));
 sky130_fd_sc_hd__a22o_1 _6471_ (.A1(\mem[21][18] ),
    .A2(_1096_),
    .B1(_1098_),
    .B2(\mem[17][18] ),
    .X(_3083_));
 sky130_fd_sc_hd__a221o_1 _6472_ (.A1(\mem[2][18] ),
    .A2(_1092_),
    .B1(_1094_),
    .B2(\mem[23][18] ),
    .C1(_3083_),
    .X(_3084_));
 sky130_fd_sc_hd__or4_4 _6473_ (.A(_3076_),
    .B(_3080_),
    .C(_3082_),
    .D(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__clkbuf_4 _6474_ (.A(_3085_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 _6475_ (.A(net18),
    .X(_3086_));
 sky130_fd_sc_hd__nand2_1 _6476_ (.A(net17),
    .B(net12),
    .Y(_3087_));
 sky130_fd_sc_hd__nand2_1 _6477_ (.A(net14),
    .B(net13),
    .Y(_3088_));
 sky130_fd_sc_hd__nand2_1 _6478_ (.A(net16),
    .B(net15),
    .Y(_3089_));
 sky130_fd_sc_hd__or3_4 _6479_ (.A(_3087_),
    .B(_3088_),
    .C(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__buf_6 _6480_ (.A(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__mux2_1 _6481_ (.A0(_3086_),
    .A1(\mem[31][0] ),
    .S(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__clkbuf_1 _6482_ (.A(_3092_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_2 _6483_ (.A(net29),
    .X(_3093_));
 sky130_fd_sc_hd__mux2_1 _6484_ (.A0(_3093_),
    .A1(\mem[31][1] ),
    .S(_3091_),
    .X(_3094_));
 sky130_fd_sc_hd__clkbuf_1 _6485_ (.A(_3094_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_2 _6486_ (.A(net40),
    .X(_3095_));
 sky130_fd_sc_hd__mux2_1 _6487_ (.A0(_3095_),
    .A1(\mem[31][2] ),
    .S(_3091_),
    .X(_3096_));
 sky130_fd_sc_hd__clkbuf_1 _6488_ (.A(_3096_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _6489_ (.A(net43),
    .X(_3097_));
 sky130_fd_sc_hd__mux2_1 _6490_ (.A0(_3097_),
    .A1(\mem[31][3] ),
    .S(_3091_),
    .X(_3098_));
 sky130_fd_sc_hd__clkbuf_1 _6491_ (.A(_3098_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_2 _6492_ (.A(net44),
    .X(_3099_));
 sky130_fd_sc_hd__mux2_1 _6493_ (.A0(_3099_),
    .A1(\mem[31][4] ),
    .S(_3091_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_1 _6494_ (.A(_3100_),
    .X(_0004_));
 sky130_fd_sc_hd__buf_2 _6495_ (.A(net45),
    .X(_3101_));
 sky130_fd_sc_hd__mux2_1 _6496_ (.A0(_3101_),
    .A1(\mem[31][5] ),
    .S(_3091_),
    .X(_3102_));
 sky130_fd_sc_hd__clkbuf_1 _6497_ (.A(_3102_),
    .X(_0005_));
 sky130_fd_sc_hd__buf_2 _6498_ (.A(net46),
    .X(_3103_));
 sky130_fd_sc_hd__mux2_1 _6499_ (.A0(_3103_),
    .A1(\mem[31][6] ),
    .S(_3091_),
    .X(_3104_));
 sky130_fd_sc_hd__clkbuf_1 _6500_ (.A(_3104_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_2 _6501_ (.A(net47),
    .X(_3105_));
 sky130_fd_sc_hd__mux2_1 _6502_ (.A0(_3105_),
    .A1(\mem[31][7] ),
    .S(_3091_),
    .X(_3106_));
 sky130_fd_sc_hd__clkbuf_1 _6503_ (.A(_3106_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_2 _6504_ (.A(net48),
    .X(_3107_));
 sky130_fd_sc_hd__mux2_1 _6505_ (.A0(_3107_),
    .A1(\mem[31][8] ),
    .S(_3091_),
    .X(_3108_));
 sky130_fd_sc_hd__clkbuf_1 _6506_ (.A(_3108_),
    .X(_0008_));
 sky130_fd_sc_hd__buf_2 _6507_ (.A(net49),
    .X(_3109_));
 sky130_fd_sc_hd__mux2_1 _6508_ (.A0(_3109_),
    .A1(\mem[31][9] ),
    .S(_3091_),
    .X(_3110_));
 sky130_fd_sc_hd__clkbuf_1 _6509_ (.A(_3110_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _6510_ (.A(net19),
    .X(_3111_));
 sky130_fd_sc_hd__buf_6 _6511_ (.A(_3090_),
    .X(_3112_));
 sky130_fd_sc_hd__mux2_1 _6512_ (.A0(_3111_),
    .A1(\mem[31][10] ),
    .S(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__clkbuf_1 _6513_ (.A(_3113_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _6514_ (.A(net20),
    .X(_3114_));
 sky130_fd_sc_hd__mux2_1 _6515_ (.A0(_3114_),
    .A1(\mem[31][11] ),
    .S(_3112_),
    .X(_3115_));
 sky130_fd_sc_hd__clkbuf_1 _6516_ (.A(_3115_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_2 _6517_ (.A(net21),
    .X(_3116_));
 sky130_fd_sc_hd__mux2_1 _6518_ (.A0(_3116_),
    .A1(\mem[31][12] ),
    .S(_3112_),
    .X(_3117_));
 sky130_fd_sc_hd__clkbuf_1 _6519_ (.A(_3117_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_2 _6520_ (.A(net22),
    .X(_3118_));
 sky130_fd_sc_hd__mux2_1 _6521_ (.A0(_3118_),
    .A1(\mem[31][13] ),
    .S(_3112_),
    .X(_3119_));
 sky130_fd_sc_hd__clkbuf_1 _6522_ (.A(_3119_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_2 _6523_ (.A(net23),
    .X(_3120_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(_3120_),
    .A1(\mem[31][14] ),
    .S(_3112_),
    .X(_3121_));
 sky130_fd_sc_hd__clkbuf_1 _6525_ (.A(_3121_),
    .X(_0014_));
 sky130_fd_sc_hd__buf_2 _6526_ (.A(net24),
    .X(_3122_));
 sky130_fd_sc_hd__mux2_1 _6527_ (.A0(_3122_),
    .A1(\mem[31][15] ),
    .S(_3112_),
    .X(_3123_));
 sky130_fd_sc_hd__clkbuf_1 _6528_ (.A(_3123_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_2 _6529_ (.A(net25),
    .X(_3124_));
 sky130_fd_sc_hd__mux2_1 _6530_ (.A0(_3124_),
    .A1(\mem[31][16] ),
    .S(_3112_),
    .X(_3125_));
 sky130_fd_sc_hd__clkbuf_1 _6531_ (.A(_3125_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_2 _6532_ (.A(net26),
    .X(_3126_));
 sky130_fd_sc_hd__mux2_1 _6533_ (.A0(_3126_),
    .A1(\mem[31][17] ),
    .S(_3112_),
    .X(_3127_));
 sky130_fd_sc_hd__clkbuf_1 _6534_ (.A(_3127_),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _6535_ (.A(net27),
    .X(_3128_));
 sky130_fd_sc_hd__mux2_1 _6536_ (.A0(_3128_),
    .A1(\mem[31][18] ),
    .S(_3112_),
    .X(_3129_));
 sky130_fd_sc_hd__clkbuf_1 _6537_ (.A(_3129_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_2 _6538_ (.A(net28),
    .X(_3130_));
 sky130_fd_sc_hd__mux2_1 _6539_ (.A0(_3130_),
    .A1(\mem[31][19] ),
    .S(_3112_),
    .X(_3131_));
 sky130_fd_sc_hd__clkbuf_1 _6540_ (.A(_3131_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _6541_ (.A(net30),
    .X(_3132_));
 sky130_fd_sc_hd__buf_4 _6542_ (.A(_3090_),
    .X(_3133_));
 sky130_fd_sc_hd__mux2_1 _6543_ (.A0(_3132_),
    .A1(\mem[31][20] ),
    .S(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__clkbuf_1 _6544_ (.A(_3134_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_2 _6545_ (.A(net31),
    .X(_3135_));
 sky130_fd_sc_hd__mux2_1 _6546_ (.A0(_3135_),
    .A1(\mem[31][21] ),
    .S(_3133_),
    .X(_3136_));
 sky130_fd_sc_hd__clkbuf_1 _6547_ (.A(_3136_),
    .X(_0021_));
 sky130_fd_sc_hd__buf_2 _6548_ (.A(net32),
    .X(_3137_));
 sky130_fd_sc_hd__mux2_1 _6549_ (.A0(_3137_),
    .A1(\mem[31][22] ),
    .S(_3133_),
    .X(_3138_));
 sky130_fd_sc_hd__clkbuf_1 _6550_ (.A(_3138_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_2 _6551_ (.A(net33),
    .X(_3139_));
 sky130_fd_sc_hd__mux2_1 _6552_ (.A0(_3139_),
    .A1(\mem[31][23] ),
    .S(_3133_),
    .X(_3140_));
 sky130_fd_sc_hd__clkbuf_1 _6553_ (.A(_3140_),
    .X(_0023_));
 sky130_fd_sc_hd__buf_2 _6554_ (.A(net34),
    .X(_3141_));
 sky130_fd_sc_hd__mux2_1 _6555_ (.A0(_3141_),
    .A1(\mem[31][24] ),
    .S(_3133_),
    .X(_3142_));
 sky130_fd_sc_hd__clkbuf_1 _6556_ (.A(_3142_),
    .X(_0024_));
 sky130_fd_sc_hd__buf_2 _6557_ (.A(net35),
    .X(_3143_));
 sky130_fd_sc_hd__mux2_1 _6558_ (.A0(_3143_),
    .A1(\mem[31][25] ),
    .S(_3133_),
    .X(_3144_));
 sky130_fd_sc_hd__clkbuf_1 _6559_ (.A(_3144_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_2 _6560_ (.A(net36),
    .X(_3145_));
 sky130_fd_sc_hd__mux2_1 _6561_ (.A0(_3145_),
    .A1(\mem[31][26] ),
    .S(_3133_),
    .X(_3146_));
 sky130_fd_sc_hd__clkbuf_1 _6562_ (.A(_3146_),
    .X(_0026_));
 sky130_fd_sc_hd__buf_2 _6563_ (.A(net37),
    .X(_3147_));
 sky130_fd_sc_hd__mux2_1 _6564_ (.A0(_3147_),
    .A1(\mem[31][27] ),
    .S(_3133_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_1 _6565_ (.A(_3148_),
    .X(_0027_));
 sky130_fd_sc_hd__buf_2 _6566_ (.A(net38),
    .X(_3149_));
 sky130_fd_sc_hd__mux2_1 _6567_ (.A0(_3149_),
    .A1(\mem[31][28] ),
    .S(_3133_),
    .X(_3150_));
 sky130_fd_sc_hd__clkbuf_1 _6568_ (.A(_3150_),
    .X(_0028_));
 sky130_fd_sc_hd__buf_2 _6569_ (.A(net39),
    .X(_3151_));
 sky130_fd_sc_hd__mux2_1 _6570_ (.A0(_3151_),
    .A1(\mem[31][29] ),
    .S(_3133_),
    .X(_3152_));
 sky130_fd_sc_hd__clkbuf_1 _6571_ (.A(_3152_),
    .X(_0029_));
 sky130_fd_sc_hd__buf_2 _6572_ (.A(net41),
    .X(_3153_));
 sky130_fd_sc_hd__mux2_1 _6573_ (.A0(_3153_),
    .A1(\mem[31][30] ),
    .S(_3090_),
    .X(_3154_));
 sky130_fd_sc_hd__clkbuf_1 _6574_ (.A(_3154_),
    .X(_0030_));
 sky130_fd_sc_hd__buf_2 _6575_ (.A(net42),
    .X(_3155_));
 sky130_fd_sc_hd__mux2_1 _6576_ (.A0(_3155_),
    .A1(\mem[31][31] ),
    .S(_3090_),
    .X(_3156_));
 sky130_fd_sc_hd__clkbuf_1 _6577_ (.A(_3156_),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_2 _6578_ (.A(net18),
    .X(_3157_));
 sky130_fd_sc_hd__nor2b_2 _6579_ (.A(net17),
    .B_N(net12),
    .Y(_3158_));
 sky130_fd_sc_hd__and2b_1 _6580_ (.A_N(net14),
    .B(net13),
    .X(_3159_));
 sky130_fd_sc_hd__nor2_2 _6581_ (.A(net16),
    .B(net15),
    .Y(_3160_));
 sky130_fd_sc_hd__and3_2 _6582_ (.A(_3158_),
    .B(_3159_),
    .C(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__buf_4 _6583_ (.A(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__mux2_1 _6584_ (.A0(\mem[1][0] ),
    .A1(_3157_),
    .S(_3162_),
    .X(_3163_));
 sky130_fd_sc_hd__clkbuf_1 _6585_ (.A(_3163_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_2 _6586_ (.A(net29),
    .X(_3164_));
 sky130_fd_sc_hd__mux2_1 _6587_ (.A0(\mem[1][1] ),
    .A1(_3164_),
    .S(_3162_),
    .X(_3165_));
 sky130_fd_sc_hd__clkbuf_1 _6588_ (.A(_3165_),
    .X(_0033_));
 sky130_fd_sc_hd__buf_2 _6589_ (.A(net40),
    .X(_3166_));
 sky130_fd_sc_hd__mux2_1 _6590_ (.A0(\mem[1][2] ),
    .A1(_3166_),
    .S(_3162_),
    .X(_3167_));
 sky130_fd_sc_hd__clkbuf_1 _6591_ (.A(_3167_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_4 _6592_ (.A(net43),
    .X(_3168_));
 sky130_fd_sc_hd__mux2_1 _6593_ (.A0(\mem[1][3] ),
    .A1(_3168_),
    .S(_3162_),
    .X(_3169_));
 sky130_fd_sc_hd__clkbuf_1 _6594_ (.A(_3169_),
    .X(_0035_));
 sky130_fd_sc_hd__buf_2 _6595_ (.A(net44),
    .X(_3170_));
 sky130_fd_sc_hd__mux2_1 _6596_ (.A0(\mem[1][4] ),
    .A1(_3170_),
    .S(_3162_),
    .X(_3171_));
 sky130_fd_sc_hd__clkbuf_1 _6597_ (.A(_3171_),
    .X(_0036_));
 sky130_fd_sc_hd__buf_2 _6598_ (.A(net45),
    .X(_3172_));
 sky130_fd_sc_hd__mux2_1 _6599_ (.A0(\mem[1][5] ),
    .A1(_3172_),
    .S(_3162_),
    .X(_3173_));
 sky130_fd_sc_hd__clkbuf_1 _6600_ (.A(_3173_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _6601_ (.A(net46),
    .X(_3174_));
 sky130_fd_sc_hd__mux2_1 _6602_ (.A0(\mem[1][6] ),
    .A1(_3174_),
    .S(_3162_),
    .X(_3175_));
 sky130_fd_sc_hd__clkbuf_1 _6603_ (.A(_3175_),
    .X(_0038_));
 sky130_fd_sc_hd__buf_2 _6604_ (.A(net47),
    .X(_3176_));
 sky130_fd_sc_hd__mux2_1 _6605_ (.A0(\mem[1][7] ),
    .A1(_3176_),
    .S(_3162_),
    .X(_3177_));
 sky130_fd_sc_hd__clkbuf_1 _6606_ (.A(_3177_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _6607_ (.A(net48),
    .X(_3178_));
 sky130_fd_sc_hd__mux2_1 _6608_ (.A0(\mem[1][8] ),
    .A1(_3178_),
    .S(_3162_),
    .X(_3179_));
 sky130_fd_sc_hd__clkbuf_1 _6609_ (.A(_3179_),
    .X(_0040_));
 sky130_fd_sc_hd__buf_2 _6610_ (.A(net49),
    .X(_3180_));
 sky130_fd_sc_hd__mux2_1 _6611_ (.A0(\mem[1][9] ),
    .A1(_3180_),
    .S(_3162_),
    .X(_3181_));
 sky130_fd_sc_hd__clkbuf_1 _6612_ (.A(_3181_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_2 _6613_ (.A(net19),
    .X(_3182_));
 sky130_fd_sc_hd__buf_4 _6614_ (.A(_3161_),
    .X(_3183_));
 sky130_fd_sc_hd__mux2_1 _6615_ (.A0(\mem[1][10] ),
    .A1(_3182_),
    .S(_3183_),
    .X(_3184_));
 sky130_fd_sc_hd__clkbuf_1 _6616_ (.A(_3184_),
    .X(_0042_));
 sky130_fd_sc_hd__buf_2 _6617_ (.A(net20),
    .X(_3185_));
 sky130_fd_sc_hd__mux2_1 _6618_ (.A0(\mem[1][11] ),
    .A1(_3185_),
    .S(_3183_),
    .X(_3186_));
 sky130_fd_sc_hd__clkbuf_1 _6619_ (.A(_3186_),
    .X(_0043_));
 sky130_fd_sc_hd__buf_2 _6620_ (.A(net21),
    .X(_3187_));
 sky130_fd_sc_hd__mux2_1 _6621_ (.A0(\mem[1][12] ),
    .A1(_3187_),
    .S(_3183_),
    .X(_3188_));
 sky130_fd_sc_hd__clkbuf_1 _6622_ (.A(_3188_),
    .X(_0044_));
 sky130_fd_sc_hd__buf_2 _6623_ (.A(net22),
    .X(_3189_));
 sky130_fd_sc_hd__mux2_1 _6624_ (.A0(\mem[1][13] ),
    .A1(_3189_),
    .S(_3183_),
    .X(_3190_));
 sky130_fd_sc_hd__clkbuf_1 _6625_ (.A(_3190_),
    .X(_0045_));
 sky130_fd_sc_hd__buf_2 _6626_ (.A(net23),
    .X(_3191_));
 sky130_fd_sc_hd__mux2_1 _6627_ (.A0(\mem[1][14] ),
    .A1(_3191_),
    .S(_3183_),
    .X(_3192_));
 sky130_fd_sc_hd__clkbuf_1 _6628_ (.A(_3192_),
    .X(_0046_));
 sky130_fd_sc_hd__buf_2 _6629_ (.A(net24),
    .X(_3193_));
 sky130_fd_sc_hd__mux2_1 _6630_ (.A0(\mem[1][15] ),
    .A1(_3193_),
    .S(_3183_),
    .X(_3194_));
 sky130_fd_sc_hd__clkbuf_1 _6631_ (.A(_3194_),
    .X(_0047_));
 sky130_fd_sc_hd__buf_2 _6632_ (.A(net25),
    .X(_3195_));
 sky130_fd_sc_hd__mux2_1 _6633_ (.A0(\mem[1][16] ),
    .A1(_3195_),
    .S(_3183_),
    .X(_3196_));
 sky130_fd_sc_hd__clkbuf_1 _6634_ (.A(_3196_),
    .X(_0048_));
 sky130_fd_sc_hd__buf_2 _6635_ (.A(net26),
    .X(_3197_));
 sky130_fd_sc_hd__mux2_1 _6636_ (.A0(\mem[1][17] ),
    .A1(_3197_),
    .S(_3183_),
    .X(_3198_));
 sky130_fd_sc_hd__clkbuf_1 _6637_ (.A(_3198_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_2 _6638_ (.A(net27),
    .X(_3199_));
 sky130_fd_sc_hd__mux2_1 _6639_ (.A0(\mem[1][18] ),
    .A1(_3199_),
    .S(_3183_),
    .X(_3200_));
 sky130_fd_sc_hd__clkbuf_1 _6640_ (.A(_3200_),
    .X(_0050_));
 sky130_fd_sc_hd__buf_2 _6641_ (.A(net28),
    .X(_3201_));
 sky130_fd_sc_hd__mux2_1 _6642_ (.A0(\mem[1][19] ),
    .A1(_3201_),
    .S(_3183_),
    .X(_3202_));
 sky130_fd_sc_hd__clkbuf_1 _6643_ (.A(_3202_),
    .X(_0051_));
 sky130_fd_sc_hd__buf_2 _6644_ (.A(net30),
    .X(_3203_));
 sky130_fd_sc_hd__buf_4 _6645_ (.A(_3161_),
    .X(_3204_));
 sky130_fd_sc_hd__mux2_1 _6646_ (.A0(\mem[1][20] ),
    .A1(_3203_),
    .S(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__clkbuf_1 _6647_ (.A(_3205_),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_4 _6648_ (.A(net31),
    .X(_3206_));
 sky130_fd_sc_hd__mux2_1 _6649_ (.A0(\mem[1][21] ),
    .A1(_3206_),
    .S(_3204_),
    .X(_3207_));
 sky130_fd_sc_hd__clkbuf_1 _6650_ (.A(_3207_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_2 _6651_ (.A(net32),
    .X(_3208_));
 sky130_fd_sc_hd__mux2_1 _6652_ (.A0(\mem[1][22] ),
    .A1(_3208_),
    .S(_3204_),
    .X(_3209_));
 sky130_fd_sc_hd__clkbuf_1 _6653_ (.A(_3209_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _6654_ (.A(net33),
    .X(_3210_));
 sky130_fd_sc_hd__mux2_1 _6655_ (.A0(\mem[1][23] ),
    .A1(_3210_),
    .S(_3204_),
    .X(_3211_));
 sky130_fd_sc_hd__clkbuf_1 _6656_ (.A(_3211_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_2 _6657_ (.A(net34),
    .X(_3212_));
 sky130_fd_sc_hd__mux2_1 _6658_ (.A0(\mem[1][24] ),
    .A1(_3212_),
    .S(_3204_),
    .X(_3213_));
 sky130_fd_sc_hd__clkbuf_1 _6659_ (.A(_3213_),
    .X(_0056_));
 sky130_fd_sc_hd__buf_2 _6660_ (.A(net35),
    .X(_3214_));
 sky130_fd_sc_hd__mux2_1 _6661_ (.A0(\mem[1][25] ),
    .A1(_3214_),
    .S(_3204_),
    .X(_3215_));
 sky130_fd_sc_hd__clkbuf_1 _6662_ (.A(_3215_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_2 _6663_ (.A(net36),
    .X(_3216_));
 sky130_fd_sc_hd__mux2_1 _6664_ (.A0(\mem[1][26] ),
    .A1(_3216_),
    .S(_3204_),
    .X(_3217_));
 sky130_fd_sc_hd__clkbuf_1 _6665_ (.A(_3217_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_2 _6666_ (.A(net37),
    .X(_3218_));
 sky130_fd_sc_hd__mux2_1 _6667_ (.A0(\mem[1][27] ),
    .A1(_3218_),
    .S(_3204_),
    .X(_3219_));
 sky130_fd_sc_hd__clkbuf_1 _6668_ (.A(_3219_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_2 _6669_ (.A(net38),
    .X(_3220_));
 sky130_fd_sc_hd__mux2_1 _6670_ (.A0(\mem[1][28] ),
    .A1(_3220_),
    .S(_3204_),
    .X(_3221_));
 sky130_fd_sc_hd__clkbuf_1 _6671_ (.A(_3221_),
    .X(_0060_));
 sky130_fd_sc_hd__buf_2 _6672_ (.A(net39),
    .X(_3222_));
 sky130_fd_sc_hd__mux2_1 _6673_ (.A0(\mem[1][29] ),
    .A1(_3222_),
    .S(_3204_),
    .X(_3223_));
 sky130_fd_sc_hd__clkbuf_1 _6674_ (.A(_3223_),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_4 _6675_ (.A(net41),
    .X(_3224_));
 sky130_fd_sc_hd__mux2_1 _6676_ (.A0(\mem[1][30] ),
    .A1(_3224_),
    .S(_3161_),
    .X(_3225_));
 sky130_fd_sc_hd__clkbuf_1 _6677_ (.A(_3225_),
    .X(_0062_));
 sky130_fd_sc_hd__buf_2 _6678_ (.A(net42),
    .X(_3226_));
 sky130_fd_sc_hd__mux2_1 _6679_ (.A0(\mem[1][31] ),
    .A1(_3226_),
    .S(_3161_),
    .X(_3227_));
 sky130_fd_sc_hd__clkbuf_1 _6680_ (.A(_3227_),
    .X(_0063_));
 sky130_fd_sc_hd__and2b_1 _6681_ (.A_N(net13),
    .B(net14),
    .X(_3228_));
 sky130_fd_sc_hd__and3_4 _6682_ (.A(_3158_),
    .B(_3160_),
    .C(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__buf_6 _6683_ (.A(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__mux2_1 _6684_ (.A0(\mem[2][0] ),
    .A1(_3157_),
    .S(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__clkbuf_1 _6685_ (.A(_3231_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _6686_ (.A0(\mem[2][1] ),
    .A1(_3164_),
    .S(_3230_),
    .X(_3232_));
 sky130_fd_sc_hd__clkbuf_1 _6687_ (.A(_3232_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _6688_ (.A0(\mem[2][2] ),
    .A1(_3166_),
    .S(_3230_),
    .X(_3233_));
 sky130_fd_sc_hd__clkbuf_1 _6689_ (.A(_3233_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _6690_ (.A0(\mem[2][3] ),
    .A1(_3168_),
    .S(_3230_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_1 _6691_ (.A(_3234_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _6692_ (.A0(\mem[2][4] ),
    .A1(_3170_),
    .S(_3230_),
    .X(_3235_));
 sky130_fd_sc_hd__clkbuf_1 _6693_ (.A(_3235_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _6694_ (.A0(\mem[2][5] ),
    .A1(_3172_),
    .S(_3230_),
    .X(_3236_));
 sky130_fd_sc_hd__clkbuf_1 _6695_ (.A(_3236_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _6696_ (.A0(\mem[2][6] ),
    .A1(_3174_),
    .S(_3230_),
    .X(_3237_));
 sky130_fd_sc_hd__clkbuf_1 _6697_ (.A(_3237_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _6698_ (.A0(\mem[2][7] ),
    .A1(_3176_),
    .S(_3230_),
    .X(_3238_));
 sky130_fd_sc_hd__clkbuf_1 _6699_ (.A(_3238_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _6700_ (.A0(\mem[2][8] ),
    .A1(_3178_),
    .S(_3230_),
    .X(_3239_));
 sky130_fd_sc_hd__clkbuf_1 _6701_ (.A(_3239_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _6702_ (.A0(\mem[2][9] ),
    .A1(_3180_),
    .S(_3230_),
    .X(_3240_));
 sky130_fd_sc_hd__clkbuf_1 _6703_ (.A(_3240_),
    .X(_0073_));
 sky130_fd_sc_hd__buf_6 _6704_ (.A(_3229_),
    .X(_3241_));
 sky130_fd_sc_hd__mux2_1 _6705_ (.A0(\mem[2][10] ),
    .A1(_3182_),
    .S(_3241_),
    .X(_3242_));
 sky130_fd_sc_hd__clkbuf_1 _6706_ (.A(_3242_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _6707_ (.A0(\mem[2][11] ),
    .A1(_3185_),
    .S(_3241_),
    .X(_3243_));
 sky130_fd_sc_hd__clkbuf_1 _6708_ (.A(_3243_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _6709_ (.A0(\mem[2][12] ),
    .A1(_3187_),
    .S(_3241_),
    .X(_3244_));
 sky130_fd_sc_hd__clkbuf_1 _6710_ (.A(_3244_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _6711_ (.A0(\mem[2][13] ),
    .A1(_3189_),
    .S(_3241_),
    .X(_3245_));
 sky130_fd_sc_hd__clkbuf_1 _6712_ (.A(_3245_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _6713_ (.A0(\mem[2][14] ),
    .A1(_3191_),
    .S(_3241_),
    .X(_3246_));
 sky130_fd_sc_hd__clkbuf_1 _6714_ (.A(_3246_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _6715_ (.A0(\mem[2][15] ),
    .A1(_3193_),
    .S(_3241_),
    .X(_3247_));
 sky130_fd_sc_hd__clkbuf_1 _6716_ (.A(_3247_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _6717_ (.A0(\mem[2][16] ),
    .A1(_3195_),
    .S(_3241_),
    .X(_3248_));
 sky130_fd_sc_hd__clkbuf_1 _6718_ (.A(_3248_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _6719_ (.A0(\mem[2][17] ),
    .A1(_3197_),
    .S(_3241_),
    .X(_3249_));
 sky130_fd_sc_hd__clkbuf_1 _6720_ (.A(_3249_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _6721_ (.A0(\mem[2][18] ),
    .A1(_3199_),
    .S(_3241_),
    .X(_3250_));
 sky130_fd_sc_hd__clkbuf_1 _6722_ (.A(_3250_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _6723_ (.A0(\mem[2][19] ),
    .A1(_3201_),
    .S(_3241_),
    .X(_3251_));
 sky130_fd_sc_hd__clkbuf_1 _6724_ (.A(_3251_),
    .X(_0083_));
 sky130_fd_sc_hd__buf_4 _6725_ (.A(_3229_),
    .X(_3252_));
 sky130_fd_sc_hd__mux2_1 _6726_ (.A0(\mem[2][20] ),
    .A1(_3203_),
    .S(_3252_),
    .X(_3253_));
 sky130_fd_sc_hd__clkbuf_1 _6727_ (.A(_3253_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _6728_ (.A0(\mem[2][21] ),
    .A1(_3206_),
    .S(_3252_),
    .X(_3254_));
 sky130_fd_sc_hd__clkbuf_1 _6729_ (.A(_3254_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _6730_ (.A0(\mem[2][22] ),
    .A1(_3208_),
    .S(_3252_),
    .X(_3255_));
 sky130_fd_sc_hd__clkbuf_1 _6731_ (.A(_3255_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _6732_ (.A0(\mem[2][23] ),
    .A1(_3210_),
    .S(_3252_),
    .X(_3256_));
 sky130_fd_sc_hd__clkbuf_1 _6733_ (.A(_3256_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _6734_ (.A0(\mem[2][24] ),
    .A1(_3212_),
    .S(_3252_),
    .X(_3257_));
 sky130_fd_sc_hd__clkbuf_1 _6735_ (.A(_3257_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _6736_ (.A0(\mem[2][25] ),
    .A1(_3214_),
    .S(_3252_),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_1 _6737_ (.A(_3258_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _6738_ (.A0(\mem[2][26] ),
    .A1(_3216_),
    .S(_3252_),
    .X(_3259_));
 sky130_fd_sc_hd__clkbuf_1 _6739_ (.A(_3259_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _6740_ (.A0(\mem[2][27] ),
    .A1(_3218_),
    .S(_3252_),
    .X(_3260_));
 sky130_fd_sc_hd__clkbuf_1 _6741_ (.A(_3260_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _6742_ (.A0(\mem[2][28] ),
    .A1(_3220_),
    .S(_3252_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_1 _6743_ (.A(_3261_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _6744_ (.A0(\mem[2][29] ),
    .A1(_3222_),
    .S(_3252_),
    .X(_3262_));
 sky130_fd_sc_hd__clkbuf_1 _6745_ (.A(_3262_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _6746_ (.A0(\mem[2][30] ),
    .A1(_3224_),
    .S(_3229_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_1 _6747_ (.A(_3263_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _6748_ (.A0(\mem[2][31] ),
    .A1(_3226_),
    .S(_3229_),
    .X(_3264_));
 sky130_fd_sc_hd__clkbuf_1 _6749_ (.A(_3264_),
    .X(_0095_));
 sky130_fd_sc_hd__and3b_1 _6750_ (.A_N(_3088_),
    .B(_3158_),
    .C(_3160_),
    .X(_3265_));
 sky130_fd_sc_hd__buf_2 _6751_ (.A(_3265_),
    .X(_3266_));
 sky130_fd_sc_hd__buf_4 _6752_ (.A(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__mux2_1 _6753_ (.A0(\mem[3][0] ),
    .A1(_3157_),
    .S(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__clkbuf_1 _6754_ (.A(_3268_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _6755_ (.A0(\mem[3][1] ),
    .A1(_3164_),
    .S(_3267_),
    .X(_3269_));
 sky130_fd_sc_hd__clkbuf_1 _6756_ (.A(_3269_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _6757_ (.A0(\mem[3][2] ),
    .A1(_3166_),
    .S(_3267_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_1 _6758_ (.A(_3270_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _6759_ (.A0(\mem[3][3] ),
    .A1(_3168_),
    .S(_3267_),
    .X(_3271_));
 sky130_fd_sc_hd__clkbuf_1 _6760_ (.A(_3271_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _6761_ (.A0(\mem[3][4] ),
    .A1(_3170_),
    .S(_3267_),
    .X(_3272_));
 sky130_fd_sc_hd__clkbuf_1 _6762_ (.A(_3272_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _6763_ (.A0(\mem[3][5] ),
    .A1(_3172_),
    .S(_3267_),
    .X(_3273_));
 sky130_fd_sc_hd__clkbuf_1 _6764_ (.A(_3273_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _6765_ (.A0(\mem[3][6] ),
    .A1(_3174_),
    .S(_3267_),
    .X(_3274_));
 sky130_fd_sc_hd__clkbuf_1 _6766_ (.A(_3274_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _6767_ (.A0(\mem[3][7] ),
    .A1(_3176_),
    .S(_3267_),
    .X(_3275_));
 sky130_fd_sc_hd__clkbuf_1 _6768_ (.A(_3275_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _6769_ (.A0(\mem[3][8] ),
    .A1(_3178_),
    .S(_3267_),
    .X(_3276_));
 sky130_fd_sc_hd__clkbuf_1 _6770_ (.A(_3276_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _6771_ (.A0(\mem[3][9] ),
    .A1(_3180_),
    .S(_3267_),
    .X(_3277_));
 sky130_fd_sc_hd__clkbuf_1 _6772_ (.A(_3277_),
    .X(_0105_));
 sky130_fd_sc_hd__buf_4 _6773_ (.A(_3266_),
    .X(_3278_));
 sky130_fd_sc_hd__mux2_1 _6774_ (.A0(\mem[3][10] ),
    .A1(_3182_),
    .S(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__clkbuf_1 _6775_ (.A(_3279_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _6776_ (.A0(\mem[3][11] ),
    .A1(_3185_),
    .S(_3278_),
    .X(_3280_));
 sky130_fd_sc_hd__clkbuf_1 _6777_ (.A(_3280_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _6778_ (.A0(\mem[3][12] ),
    .A1(_3187_),
    .S(_3278_),
    .X(_3281_));
 sky130_fd_sc_hd__clkbuf_1 _6779_ (.A(_3281_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _6780_ (.A0(\mem[3][13] ),
    .A1(_3189_),
    .S(_3278_),
    .X(_3282_));
 sky130_fd_sc_hd__clkbuf_1 _6781_ (.A(_3282_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _6782_ (.A0(\mem[3][14] ),
    .A1(_3191_),
    .S(_3278_),
    .X(_3283_));
 sky130_fd_sc_hd__clkbuf_1 _6783_ (.A(_3283_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _6784_ (.A0(\mem[3][15] ),
    .A1(_3193_),
    .S(_3278_),
    .X(_3284_));
 sky130_fd_sc_hd__clkbuf_1 _6785_ (.A(_3284_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _6786_ (.A0(\mem[3][16] ),
    .A1(_3195_),
    .S(_3278_),
    .X(_3285_));
 sky130_fd_sc_hd__clkbuf_1 _6787_ (.A(_3285_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _6788_ (.A0(\mem[3][17] ),
    .A1(_3197_),
    .S(_3278_),
    .X(_3286_));
 sky130_fd_sc_hd__clkbuf_1 _6789_ (.A(_3286_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _6790_ (.A0(\mem[3][18] ),
    .A1(_3199_),
    .S(_3278_),
    .X(_3287_));
 sky130_fd_sc_hd__clkbuf_1 _6791_ (.A(_3287_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _6792_ (.A0(\mem[3][19] ),
    .A1(_3201_),
    .S(_3278_),
    .X(_3288_));
 sky130_fd_sc_hd__clkbuf_1 _6793_ (.A(_3288_),
    .X(_0115_));
 sky130_fd_sc_hd__buf_4 _6794_ (.A(_3266_),
    .X(_3289_));
 sky130_fd_sc_hd__mux2_1 _6795_ (.A0(\mem[3][20] ),
    .A1(_3203_),
    .S(_3289_),
    .X(_3290_));
 sky130_fd_sc_hd__clkbuf_1 _6796_ (.A(_3290_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _6797_ (.A0(\mem[3][21] ),
    .A1(_3206_),
    .S(_3289_),
    .X(_3291_));
 sky130_fd_sc_hd__clkbuf_1 _6798_ (.A(_3291_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _6799_ (.A0(\mem[3][22] ),
    .A1(_3208_),
    .S(_3289_),
    .X(_3292_));
 sky130_fd_sc_hd__clkbuf_1 _6800_ (.A(_3292_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _6801_ (.A0(\mem[3][23] ),
    .A1(_3210_),
    .S(_3289_),
    .X(_3293_));
 sky130_fd_sc_hd__clkbuf_1 _6802_ (.A(_3293_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _6803_ (.A0(\mem[3][24] ),
    .A1(_3212_),
    .S(_3289_),
    .X(_3294_));
 sky130_fd_sc_hd__clkbuf_1 _6804_ (.A(_3294_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _6805_ (.A0(\mem[3][25] ),
    .A1(_3214_),
    .S(_3289_),
    .X(_3295_));
 sky130_fd_sc_hd__clkbuf_1 _6806_ (.A(_3295_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _6807_ (.A0(\mem[3][26] ),
    .A1(_3216_),
    .S(_3289_),
    .X(_3296_));
 sky130_fd_sc_hd__clkbuf_1 _6808_ (.A(_3296_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _6809_ (.A0(\mem[3][27] ),
    .A1(_3218_),
    .S(_3289_),
    .X(_3297_));
 sky130_fd_sc_hd__clkbuf_1 _6810_ (.A(_3297_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _6811_ (.A0(\mem[3][28] ),
    .A1(_3220_),
    .S(_3289_),
    .X(_3298_));
 sky130_fd_sc_hd__clkbuf_1 _6812_ (.A(_3298_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _6813_ (.A0(\mem[3][29] ),
    .A1(_3222_),
    .S(_3289_),
    .X(_3299_));
 sky130_fd_sc_hd__clkbuf_1 _6814_ (.A(_3299_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _6815_ (.A0(\mem[3][30] ),
    .A1(_3224_),
    .S(_3266_),
    .X(_3300_));
 sky130_fd_sc_hd__clkbuf_1 _6816_ (.A(_3300_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _6817_ (.A0(\mem[3][31] ),
    .A1(_3226_),
    .S(_3266_),
    .X(_3301_));
 sky130_fd_sc_hd__clkbuf_1 _6818_ (.A(_3301_),
    .X(_0127_));
 sky130_fd_sc_hd__nor2_2 _6819_ (.A(net14),
    .B(net13),
    .Y(_3302_));
 sky130_fd_sc_hd__and2b_1 _6820_ (.A_N(net16),
    .B(net15),
    .X(_3303_));
 sky130_fd_sc_hd__and3_4 _6821_ (.A(_3158_),
    .B(_3302_),
    .C(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__buf_6 _6822_ (.A(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__mux2_1 _6823_ (.A0(\mem[4][0] ),
    .A1(_3157_),
    .S(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__clkbuf_1 _6824_ (.A(_3306_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _6825_ (.A0(\mem[4][1] ),
    .A1(_3164_),
    .S(_3305_),
    .X(_3307_));
 sky130_fd_sc_hd__clkbuf_1 _6826_ (.A(_3307_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _6827_ (.A0(\mem[4][2] ),
    .A1(_3166_),
    .S(_3305_),
    .X(_3308_));
 sky130_fd_sc_hd__clkbuf_1 _6828_ (.A(_3308_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _6829_ (.A0(\mem[4][3] ),
    .A1(_3168_),
    .S(_3305_),
    .X(_3309_));
 sky130_fd_sc_hd__clkbuf_1 _6830_ (.A(_3309_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _6831_ (.A0(\mem[4][4] ),
    .A1(_3170_),
    .S(_3305_),
    .X(_3310_));
 sky130_fd_sc_hd__clkbuf_1 _6832_ (.A(_3310_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _6833_ (.A0(\mem[4][5] ),
    .A1(_3172_),
    .S(_3305_),
    .X(_3311_));
 sky130_fd_sc_hd__clkbuf_1 _6834_ (.A(_3311_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _6835_ (.A0(\mem[4][6] ),
    .A1(_3174_),
    .S(_3305_),
    .X(_3312_));
 sky130_fd_sc_hd__clkbuf_1 _6836_ (.A(_3312_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _6837_ (.A0(\mem[4][7] ),
    .A1(_3176_),
    .S(_3305_),
    .X(_3313_));
 sky130_fd_sc_hd__clkbuf_1 _6838_ (.A(_3313_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _6839_ (.A0(\mem[4][8] ),
    .A1(_3178_),
    .S(_3305_),
    .X(_3314_));
 sky130_fd_sc_hd__clkbuf_1 _6840_ (.A(_3314_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _6841_ (.A0(\mem[4][9] ),
    .A1(_3180_),
    .S(_3305_),
    .X(_3315_));
 sky130_fd_sc_hd__clkbuf_1 _6842_ (.A(_3315_),
    .X(_0137_));
 sky130_fd_sc_hd__buf_6 _6843_ (.A(_3304_),
    .X(_3316_));
 sky130_fd_sc_hd__mux2_1 _6844_ (.A0(\mem[4][10] ),
    .A1(_3182_),
    .S(_3316_),
    .X(_3317_));
 sky130_fd_sc_hd__clkbuf_1 _6845_ (.A(_3317_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _6846_ (.A0(\mem[4][11] ),
    .A1(_3185_),
    .S(_3316_),
    .X(_3318_));
 sky130_fd_sc_hd__clkbuf_1 _6847_ (.A(_3318_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _6848_ (.A0(\mem[4][12] ),
    .A1(_3187_),
    .S(_3316_),
    .X(_3319_));
 sky130_fd_sc_hd__clkbuf_1 _6849_ (.A(_3319_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _6850_ (.A0(\mem[4][13] ),
    .A1(_3189_),
    .S(_3316_),
    .X(_3320_));
 sky130_fd_sc_hd__clkbuf_1 _6851_ (.A(_3320_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _6852_ (.A0(\mem[4][14] ),
    .A1(_3191_),
    .S(_3316_),
    .X(_3321_));
 sky130_fd_sc_hd__clkbuf_1 _6853_ (.A(_3321_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _6854_ (.A0(\mem[4][15] ),
    .A1(_3193_),
    .S(_3316_),
    .X(_3322_));
 sky130_fd_sc_hd__clkbuf_1 _6855_ (.A(_3322_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _6856_ (.A0(\mem[4][16] ),
    .A1(_3195_),
    .S(_3316_),
    .X(_3323_));
 sky130_fd_sc_hd__clkbuf_1 _6857_ (.A(_3323_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _6858_ (.A0(\mem[4][17] ),
    .A1(_3197_),
    .S(_3316_),
    .X(_3324_));
 sky130_fd_sc_hd__clkbuf_1 _6859_ (.A(_3324_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _6860_ (.A0(\mem[4][18] ),
    .A1(_3199_),
    .S(_3316_),
    .X(_3325_));
 sky130_fd_sc_hd__clkbuf_1 _6861_ (.A(_3325_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _6862_ (.A0(\mem[4][19] ),
    .A1(_3201_),
    .S(_3316_),
    .X(_3326_));
 sky130_fd_sc_hd__clkbuf_1 _6863_ (.A(_3326_),
    .X(_0147_));
 sky130_fd_sc_hd__buf_4 _6864_ (.A(_3304_),
    .X(_3327_));
 sky130_fd_sc_hd__mux2_1 _6865_ (.A0(\mem[4][20] ),
    .A1(_3203_),
    .S(_3327_),
    .X(_3328_));
 sky130_fd_sc_hd__clkbuf_1 _6866_ (.A(_3328_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _6867_ (.A0(\mem[4][21] ),
    .A1(_3206_),
    .S(_3327_),
    .X(_3329_));
 sky130_fd_sc_hd__clkbuf_1 _6868_ (.A(_3329_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _6869_ (.A0(\mem[4][22] ),
    .A1(_3208_),
    .S(_3327_),
    .X(_3330_));
 sky130_fd_sc_hd__clkbuf_1 _6870_ (.A(_3330_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _6871_ (.A0(\mem[4][23] ),
    .A1(_3210_),
    .S(_3327_),
    .X(_3331_));
 sky130_fd_sc_hd__clkbuf_1 _6872_ (.A(_3331_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _6873_ (.A0(\mem[4][24] ),
    .A1(_3212_),
    .S(_3327_),
    .X(_3332_));
 sky130_fd_sc_hd__clkbuf_1 _6874_ (.A(_3332_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _6875_ (.A0(\mem[4][25] ),
    .A1(_3214_),
    .S(_3327_),
    .X(_3333_));
 sky130_fd_sc_hd__clkbuf_1 _6876_ (.A(_3333_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _6877_ (.A0(\mem[4][26] ),
    .A1(_3216_),
    .S(_3327_),
    .X(_3334_));
 sky130_fd_sc_hd__clkbuf_1 _6878_ (.A(_3334_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _6879_ (.A0(\mem[4][27] ),
    .A1(_3218_),
    .S(_3327_),
    .X(_3335_));
 sky130_fd_sc_hd__clkbuf_1 _6880_ (.A(_3335_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _6881_ (.A0(\mem[4][28] ),
    .A1(_3220_),
    .S(_3327_),
    .X(_3336_));
 sky130_fd_sc_hd__clkbuf_1 _6882_ (.A(_3336_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _6883_ (.A0(\mem[4][29] ),
    .A1(_3222_),
    .S(_3327_),
    .X(_3337_));
 sky130_fd_sc_hd__clkbuf_1 _6884_ (.A(_3337_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _6885_ (.A0(\mem[4][30] ),
    .A1(_3224_),
    .S(_3304_),
    .X(_3338_));
 sky130_fd_sc_hd__clkbuf_1 _6886_ (.A(_3338_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _6887_ (.A0(\mem[4][31] ),
    .A1(_3226_),
    .S(_3304_),
    .X(_3339_));
 sky130_fd_sc_hd__clkbuf_1 _6888_ (.A(_3339_),
    .X(_0159_));
 sky130_fd_sc_hd__or2b_1 _6889_ (.A(net14),
    .B_N(net13),
    .X(_3340_));
 sky130_fd_sc_hd__or2b_1 _6890_ (.A(net16),
    .B_N(net15),
    .X(_3341_));
 sky130_fd_sc_hd__a21bo_1 _6891_ (.A1(_3160_),
    .A2(_3302_),
    .B1_N(_3158_),
    .X(_3342_));
 sky130_fd_sc_hd__or3_4 _6892_ (.A(_3340_),
    .B(_3341_),
    .C(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__buf_4 _6893_ (.A(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__mux2_1 _6894_ (.A0(_3086_),
    .A1(\mem[5][0] ),
    .S(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__clkbuf_1 _6895_ (.A(_3345_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _6896_ (.A0(_3093_),
    .A1(\mem[5][1] ),
    .S(_3344_),
    .X(_3346_));
 sky130_fd_sc_hd__clkbuf_1 _6897_ (.A(_3346_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _6898_ (.A0(_3095_),
    .A1(\mem[5][2] ),
    .S(_3344_),
    .X(_3347_));
 sky130_fd_sc_hd__clkbuf_1 _6899_ (.A(_3347_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _6900_ (.A0(_3097_),
    .A1(\mem[5][3] ),
    .S(_3344_),
    .X(_3348_));
 sky130_fd_sc_hd__clkbuf_1 _6901_ (.A(_3348_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _6902_ (.A0(_3099_),
    .A1(\mem[5][4] ),
    .S(_3344_),
    .X(_3349_));
 sky130_fd_sc_hd__clkbuf_1 _6903_ (.A(_3349_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _6904_ (.A0(_3101_),
    .A1(\mem[5][5] ),
    .S(_3344_),
    .X(_3350_));
 sky130_fd_sc_hd__clkbuf_1 _6905_ (.A(_3350_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _6906_ (.A0(_3103_),
    .A1(\mem[5][6] ),
    .S(_3344_),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_1 _6907_ (.A(_3351_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _6908_ (.A0(_3105_),
    .A1(\mem[5][7] ),
    .S(_3344_),
    .X(_3352_));
 sky130_fd_sc_hd__clkbuf_1 _6909_ (.A(_3352_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _6910_ (.A0(_3107_),
    .A1(\mem[5][8] ),
    .S(_3344_),
    .X(_3353_));
 sky130_fd_sc_hd__clkbuf_1 _6911_ (.A(_3353_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _6912_ (.A0(_3109_),
    .A1(\mem[5][9] ),
    .S(_3344_),
    .X(_3354_));
 sky130_fd_sc_hd__clkbuf_1 _6913_ (.A(_3354_),
    .X(_0169_));
 sky130_fd_sc_hd__buf_4 _6914_ (.A(_3343_),
    .X(_3355_));
 sky130_fd_sc_hd__mux2_1 _6915_ (.A0(_3111_),
    .A1(\mem[5][10] ),
    .S(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_1 _6916_ (.A(_3356_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _6917_ (.A0(_3114_),
    .A1(\mem[5][11] ),
    .S(_3355_),
    .X(_3357_));
 sky130_fd_sc_hd__clkbuf_1 _6918_ (.A(_3357_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _6919_ (.A0(_3116_),
    .A1(\mem[5][12] ),
    .S(_3355_),
    .X(_3358_));
 sky130_fd_sc_hd__clkbuf_1 _6920_ (.A(_3358_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _6921_ (.A0(_3118_),
    .A1(\mem[5][13] ),
    .S(_3355_),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_1 _6922_ (.A(_3359_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _6923_ (.A0(_3120_),
    .A1(\mem[5][14] ),
    .S(_3355_),
    .X(_3360_));
 sky130_fd_sc_hd__clkbuf_1 _6924_ (.A(_3360_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _6925_ (.A0(_3122_),
    .A1(\mem[5][15] ),
    .S(_3355_),
    .X(_3361_));
 sky130_fd_sc_hd__clkbuf_1 _6926_ (.A(_3361_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _6927_ (.A0(_3124_),
    .A1(\mem[5][16] ),
    .S(_3355_),
    .X(_3362_));
 sky130_fd_sc_hd__clkbuf_1 _6928_ (.A(_3362_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _6929_ (.A0(_3126_),
    .A1(\mem[5][17] ),
    .S(_3355_),
    .X(_3363_));
 sky130_fd_sc_hd__clkbuf_1 _6930_ (.A(_3363_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _6931_ (.A0(_3128_),
    .A1(\mem[5][18] ),
    .S(_3355_),
    .X(_3364_));
 sky130_fd_sc_hd__clkbuf_1 _6932_ (.A(_3364_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _6933_ (.A0(_3130_),
    .A1(\mem[5][19] ),
    .S(_3355_),
    .X(_3365_));
 sky130_fd_sc_hd__clkbuf_1 _6934_ (.A(_3365_),
    .X(_0179_));
 sky130_fd_sc_hd__buf_4 _6935_ (.A(_3343_),
    .X(_3366_));
 sky130_fd_sc_hd__mux2_1 _6936_ (.A0(_3132_),
    .A1(\mem[5][20] ),
    .S(_3366_),
    .X(_3367_));
 sky130_fd_sc_hd__clkbuf_1 _6937_ (.A(_3367_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _6938_ (.A0(_3135_),
    .A1(\mem[5][21] ),
    .S(_3366_),
    .X(_3368_));
 sky130_fd_sc_hd__clkbuf_1 _6939_ (.A(_3368_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _6940_ (.A0(_3137_),
    .A1(\mem[5][22] ),
    .S(_3366_),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_1 _6941_ (.A(_3369_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _6942_ (.A0(_3139_),
    .A1(\mem[5][23] ),
    .S(_3366_),
    .X(_3370_));
 sky130_fd_sc_hd__clkbuf_1 _6943_ (.A(_3370_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _6944_ (.A0(_3141_),
    .A1(\mem[5][24] ),
    .S(_3366_),
    .X(_3371_));
 sky130_fd_sc_hd__clkbuf_1 _6945_ (.A(_3371_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _6946_ (.A0(_3143_),
    .A1(\mem[5][25] ),
    .S(_3366_),
    .X(_3372_));
 sky130_fd_sc_hd__clkbuf_1 _6947_ (.A(_3372_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _6948_ (.A0(_3145_),
    .A1(\mem[5][26] ),
    .S(_3366_),
    .X(_3373_));
 sky130_fd_sc_hd__clkbuf_1 _6949_ (.A(_3373_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _6950_ (.A0(_3147_),
    .A1(\mem[5][27] ),
    .S(_3366_),
    .X(_3374_));
 sky130_fd_sc_hd__clkbuf_1 _6951_ (.A(_3374_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _6952_ (.A0(_3149_),
    .A1(\mem[5][28] ),
    .S(_3366_),
    .X(_3375_));
 sky130_fd_sc_hd__clkbuf_1 _6953_ (.A(_3375_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _6954_ (.A0(_3151_),
    .A1(\mem[5][29] ),
    .S(_3366_),
    .X(_3376_));
 sky130_fd_sc_hd__clkbuf_1 _6955_ (.A(_3376_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _6956_ (.A0(_3153_),
    .A1(\mem[5][30] ),
    .S(_3343_),
    .X(_3377_));
 sky130_fd_sc_hd__clkbuf_1 _6957_ (.A(_3377_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _6958_ (.A0(_3155_),
    .A1(\mem[5][31] ),
    .S(_3343_),
    .X(_3378_));
 sky130_fd_sc_hd__clkbuf_1 _6959_ (.A(_3378_),
    .X(_0191_));
 sky130_fd_sc_hd__or2b_1 _6960_ (.A(net13),
    .B_N(net14),
    .X(_3379_));
 sky130_fd_sc_hd__or3_4 _6961_ (.A(_3379_),
    .B(_3341_),
    .C(_3342_),
    .X(_3380_));
 sky130_fd_sc_hd__buf_6 _6962_ (.A(_3380_),
    .X(_3381_));
 sky130_fd_sc_hd__mux2_1 _6963_ (.A0(_3086_),
    .A1(\mem[6][0] ),
    .S(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__clkbuf_1 _6964_ (.A(_3382_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _6965_ (.A0(_3093_),
    .A1(\mem[6][1] ),
    .S(_3381_),
    .X(_3383_));
 sky130_fd_sc_hd__clkbuf_1 _6966_ (.A(_3383_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _6967_ (.A0(_3095_),
    .A1(\mem[6][2] ),
    .S(_3381_),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_1 _6968_ (.A(_3384_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _6969_ (.A0(_3097_),
    .A1(\mem[6][3] ),
    .S(_3381_),
    .X(_3385_));
 sky130_fd_sc_hd__clkbuf_1 _6970_ (.A(_3385_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _6971_ (.A0(_3099_),
    .A1(\mem[6][4] ),
    .S(_3381_),
    .X(_3386_));
 sky130_fd_sc_hd__clkbuf_1 _6972_ (.A(_3386_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _6973_ (.A0(_3101_),
    .A1(\mem[6][5] ),
    .S(_3381_),
    .X(_3387_));
 sky130_fd_sc_hd__clkbuf_1 _6974_ (.A(_3387_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _6975_ (.A0(_3103_),
    .A1(\mem[6][6] ),
    .S(_3381_),
    .X(_3388_));
 sky130_fd_sc_hd__clkbuf_1 _6976_ (.A(_3388_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _6977_ (.A0(_3105_),
    .A1(\mem[6][7] ),
    .S(_3381_),
    .X(_3389_));
 sky130_fd_sc_hd__clkbuf_1 _6978_ (.A(_3389_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _6979_ (.A0(_3107_),
    .A1(\mem[6][8] ),
    .S(_3381_),
    .X(_3390_));
 sky130_fd_sc_hd__clkbuf_1 _6980_ (.A(_3390_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _6981_ (.A0(_3109_),
    .A1(\mem[6][9] ),
    .S(_3381_),
    .X(_3391_));
 sky130_fd_sc_hd__clkbuf_1 _6982_ (.A(_3391_),
    .X(_0201_));
 sky130_fd_sc_hd__buf_6 _6983_ (.A(_3380_),
    .X(_3392_));
 sky130_fd_sc_hd__mux2_1 _6984_ (.A0(_3111_),
    .A1(\mem[6][10] ),
    .S(_3392_),
    .X(_3393_));
 sky130_fd_sc_hd__clkbuf_1 _6985_ (.A(_3393_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _6986_ (.A0(_3114_),
    .A1(\mem[6][11] ),
    .S(_3392_),
    .X(_3394_));
 sky130_fd_sc_hd__clkbuf_1 _6987_ (.A(_3394_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _6988_ (.A0(_3116_),
    .A1(\mem[6][12] ),
    .S(_3392_),
    .X(_3395_));
 sky130_fd_sc_hd__clkbuf_1 _6989_ (.A(_3395_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _6990_ (.A0(_3118_),
    .A1(\mem[6][13] ),
    .S(_3392_),
    .X(_3396_));
 sky130_fd_sc_hd__clkbuf_1 _6991_ (.A(_3396_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _6992_ (.A0(_3120_),
    .A1(\mem[6][14] ),
    .S(_3392_),
    .X(_3397_));
 sky130_fd_sc_hd__clkbuf_1 _6993_ (.A(_3397_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _6994_ (.A0(_3122_),
    .A1(\mem[6][15] ),
    .S(_3392_),
    .X(_3398_));
 sky130_fd_sc_hd__clkbuf_1 _6995_ (.A(_3398_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _6996_ (.A0(_3124_),
    .A1(\mem[6][16] ),
    .S(_3392_),
    .X(_3399_));
 sky130_fd_sc_hd__clkbuf_1 _6997_ (.A(_3399_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _6998_ (.A0(_3126_),
    .A1(\mem[6][17] ),
    .S(_3392_),
    .X(_3400_));
 sky130_fd_sc_hd__clkbuf_1 _6999_ (.A(_3400_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _7000_ (.A0(_3128_),
    .A1(\mem[6][18] ),
    .S(_3392_),
    .X(_3401_));
 sky130_fd_sc_hd__clkbuf_1 _7001_ (.A(_3401_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _7002_ (.A0(_3130_),
    .A1(\mem[6][19] ),
    .S(_3392_),
    .X(_3402_));
 sky130_fd_sc_hd__clkbuf_1 _7003_ (.A(_3402_),
    .X(_0211_));
 sky130_fd_sc_hd__buf_4 _7004_ (.A(_3380_),
    .X(_3403_));
 sky130_fd_sc_hd__mux2_1 _7005_ (.A0(_3132_),
    .A1(\mem[6][20] ),
    .S(_3403_),
    .X(_3404_));
 sky130_fd_sc_hd__clkbuf_1 _7006_ (.A(_3404_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _7007_ (.A0(_3135_),
    .A1(\mem[6][21] ),
    .S(_3403_),
    .X(_3405_));
 sky130_fd_sc_hd__clkbuf_1 _7008_ (.A(_3405_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _7009_ (.A0(_3137_),
    .A1(\mem[6][22] ),
    .S(_3403_),
    .X(_3406_));
 sky130_fd_sc_hd__clkbuf_1 _7010_ (.A(_3406_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _7011_ (.A0(_3139_),
    .A1(\mem[6][23] ),
    .S(_3403_),
    .X(_3407_));
 sky130_fd_sc_hd__clkbuf_1 _7012_ (.A(_3407_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _7013_ (.A0(_3141_),
    .A1(\mem[6][24] ),
    .S(_3403_),
    .X(_3408_));
 sky130_fd_sc_hd__clkbuf_1 _7014_ (.A(_3408_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _7015_ (.A0(_3143_),
    .A1(\mem[6][25] ),
    .S(_3403_),
    .X(_3409_));
 sky130_fd_sc_hd__clkbuf_1 _7016_ (.A(_3409_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _7017_ (.A0(_3145_),
    .A1(\mem[6][26] ),
    .S(_3403_),
    .X(_3410_));
 sky130_fd_sc_hd__clkbuf_1 _7018_ (.A(_3410_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _7019_ (.A0(_3147_),
    .A1(\mem[6][27] ),
    .S(_3403_),
    .X(_3411_));
 sky130_fd_sc_hd__clkbuf_1 _7020_ (.A(_3411_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _7021_ (.A0(_3149_),
    .A1(\mem[6][28] ),
    .S(_3403_),
    .X(_3412_));
 sky130_fd_sc_hd__clkbuf_1 _7022_ (.A(_3412_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _7023_ (.A0(_3151_),
    .A1(\mem[6][29] ),
    .S(_3403_),
    .X(_3413_));
 sky130_fd_sc_hd__clkbuf_1 _7024_ (.A(_3413_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _7025_ (.A0(_3153_),
    .A1(\mem[6][30] ),
    .S(_3380_),
    .X(_3414_));
 sky130_fd_sc_hd__clkbuf_1 _7026_ (.A(_3414_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _7027_ (.A0(_3155_),
    .A1(\mem[6][31] ),
    .S(_3380_),
    .X(_3415_));
 sky130_fd_sc_hd__clkbuf_1 _7028_ (.A(_3415_),
    .X(_0223_));
 sky130_fd_sc_hd__or3_4 _7029_ (.A(_3088_),
    .B(_3341_),
    .C(_3342_),
    .X(_3416_));
 sky130_fd_sc_hd__buf_6 _7030_ (.A(_3416_),
    .X(_3417_));
 sky130_fd_sc_hd__mux2_1 _7031_ (.A0(_3086_),
    .A1(\mem[7][0] ),
    .S(_3417_),
    .X(_3418_));
 sky130_fd_sc_hd__clkbuf_1 _7032_ (.A(_3418_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _7033_ (.A0(_3093_),
    .A1(\mem[7][1] ),
    .S(_3417_),
    .X(_3419_));
 sky130_fd_sc_hd__clkbuf_1 _7034_ (.A(_3419_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _7035_ (.A0(_3095_),
    .A1(\mem[7][2] ),
    .S(_3417_),
    .X(_3420_));
 sky130_fd_sc_hd__clkbuf_1 _7036_ (.A(_3420_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _7037_ (.A0(_3097_),
    .A1(\mem[7][3] ),
    .S(_3417_),
    .X(_3421_));
 sky130_fd_sc_hd__clkbuf_1 _7038_ (.A(_3421_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _7039_ (.A0(_3099_),
    .A1(\mem[7][4] ),
    .S(_3417_),
    .X(_3422_));
 sky130_fd_sc_hd__clkbuf_1 _7040_ (.A(_3422_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _7041_ (.A0(_3101_),
    .A1(\mem[7][5] ),
    .S(_3417_),
    .X(_3423_));
 sky130_fd_sc_hd__clkbuf_1 _7042_ (.A(_3423_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _7043_ (.A0(_3103_),
    .A1(\mem[7][6] ),
    .S(_3417_),
    .X(_3424_));
 sky130_fd_sc_hd__clkbuf_1 _7044_ (.A(_3424_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _7045_ (.A0(_3105_),
    .A1(\mem[7][7] ),
    .S(_3417_),
    .X(_3425_));
 sky130_fd_sc_hd__clkbuf_1 _7046_ (.A(_3425_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _7047_ (.A0(_3107_),
    .A1(\mem[7][8] ),
    .S(_3417_),
    .X(_3426_));
 sky130_fd_sc_hd__clkbuf_1 _7048_ (.A(_3426_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _7049_ (.A0(_3109_),
    .A1(\mem[7][9] ),
    .S(_3417_),
    .X(_3427_));
 sky130_fd_sc_hd__clkbuf_1 _7050_ (.A(_3427_),
    .X(_0233_));
 sky130_fd_sc_hd__buf_6 _7051_ (.A(_3416_),
    .X(_3428_));
 sky130_fd_sc_hd__mux2_1 _7052_ (.A0(_3111_),
    .A1(\mem[7][10] ),
    .S(_3428_),
    .X(_3429_));
 sky130_fd_sc_hd__clkbuf_1 _7053_ (.A(_3429_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _7054_ (.A0(_3114_),
    .A1(\mem[7][11] ),
    .S(_3428_),
    .X(_3430_));
 sky130_fd_sc_hd__clkbuf_1 _7055_ (.A(_3430_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _7056_ (.A0(_3116_),
    .A1(\mem[7][12] ),
    .S(_3428_),
    .X(_3431_));
 sky130_fd_sc_hd__clkbuf_1 _7057_ (.A(_3431_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _7058_ (.A0(_3118_),
    .A1(\mem[7][13] ),
    .S(_3428_),
    .X(_3432_));
 sky130_fd_sc_hd__clkbuf_1 _7059_ (.A(_3432_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _7060_ (.A0(_3120_),
    .A1(\mem[7][14] ),
    .S(_3428_),
    .X(_3433_));
 sky130_fd_sc_hd__clkbuf_1 _7061_ (.A(_3433_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _7062_ (.A0(_3122_),
    .A1(\mem[7][15] ),
    .S(_3428_),
    .X(_3434_));
 sky130_fd_sc_hd__clkbuf_1 _7063_ (.A(_3434_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _7064_ (.A0(_3124_),
    .A1(\mem[7][16] ),
    .S(_3428_),
    .X(_3435_));
 sky130_fd_sc_hd__clkbuf_1 _7065_ (.A(_3435_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _7066_ (.A0(_3126_),
    .A1(\mem[7][17] ),
    .S(_3428_),
    .X(_3436_));
 sky130_fd_sc_hd__clkbuf_1 _7067_ (.A(_3436_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _7068_ (.A0(_3128_),
    .A1(\mem[7][18] ),
    .S(_3428_),
    .X(_3437_));
 sky130_fd_sc_hd__clkbuf_1 _7069_ (.A(_3437_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _7070_ (.A0(_3130_),
    .A1(\mem[7][19] ),
    .S(_3428_),
    .X(_3438_));
 sky130_fd_sc_hd__clkbuf_1 _7071_ (.A(_3438_),
    .X(_0243_));
 sky130_fd_sc_hd__buf_4 _7072_ (.A(_3416_),
    .X(_3439_));
 sky130_fd_sc_hd__mux2_1 _7073_ (.A0(_3132_),
    .A1(\mem[7][20] ),
    .S(_3439_),
    .X(_3440_));
 sky130_fd_sc_hd__clkbuf_1 _7074_ (.A(_3440_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _7075_ (.A0(_3135_),
    .A1(\mem[7][21] ),
    .S(_3439_),
    .X(_3441_));
 sky130_fd_sc_hd__clkbuf_1 _7076_ (.A(_3441_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _7077_ (.A0(_3137_),
    .A1(\mem[7][22] ),
    .S(_3439_),
    .X(_3442_));
 sky130_fd_sc_hd__clkbuf_1 _7078_ (.A(_3442_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _7079_ (.A0(_3139_),
    .A1(\mem[7][23] ),
    .S(_3439_),
    .X(_3443_));
 sky130_fd_sc_hd__clkbuf_1 _7080_ (.A(_3443_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _7081_ (.A0(_3141_),
    .A1(\mem[7][24] ),
    .S(_3439_),
    .X(_3444_));
 sky130_fd_sc_hd__clkbuf_1 _7082_ (.A(_3444_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _7083_ (.A0(_3143_),
    .A1(\mem[7][25] ),
    .S(_3439_),
    .X(_3445_));
 sky130_fd_sc_hd__clkbuf_1 _7084_ (.A(_3445_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _7085_ (.A0(_3145_),
    .A1(\mem[7][26] ),
    .S(_3439_),
    .X(_3446_));
 sky130_fd_sc_hd__clkbuf_1 _7086_ (.A(_3446_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _7087_ (.A0(_3147_),
    .A1(\mem[7][27] ),
    .S(_3439_),
    .X(_3447_));
 sky130_fd_sc_hd__clkbuf_1 _7088_ (.A(_3447_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _7089_ (.A0(_3149_),
    .A1(\mem[7][28] ),
    .S(_3439_),
    .X(_3448_));
 sky130_fd_sc_hd__clkbuf_1 _7090_ (.A(_3448_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _7091_ (.A0(_3151_),
    .A1(\mem[7][29] ),
    .S(_3439_),
    .X(_3449_));
 sky130_fd_sc_hd__clkbuf_1 _7092_ (.A(_3449_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _7093_ (.A0(_3153_),
    .A1(\mem[7][30] ),
    .S(_3416_),
    .X(_3450_));
 sky130_fd_sc_hd__clkbuf_1 _7094_ (.A(_3450_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _7095_ (.A0(_3155_),
    .A1(\mem[7][31] ),
    .S(_3416_),
    .X(_3451_));
 sky130_fd_sc_hd__clkbuf_1 _7096_ (.A(_3451_),
    .X(_0255_));
 sky130_fd_sc_hd__and2b_1 _7097_ (.A_N(net15),
    .B(net16),
    .X(_3452_));
 sky130_fd_sc_hd__and3_2 _7098_ (.A(_3158_),
    .B(_3302_),
    .C(_3452_),
    .X(_3453_));
 sky130_fd_sc_hd__buf_6 _7099_ (.A(_3453_),
    .X(_3454_));
 sky130_fd_sc_hd__mux2_1 _7100_ (.A0(\mem[8][0] ),
    .A1(_3157_),
    .S(_3454_),
    .X(_3455_));
 sky130_fd_sc_hd__clkbuf_1 _7101_ (.A(_3455_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _7102_ (.A0(\mem[8][1] ),
    .A1(_3164_),
    .S(_3454_),
    .X(_3456_));
 sky130_fd_sc_hd__clkbuf_1 _7103_ (.A(_3456_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _7104_ (.A0(\mem[8][2] ),
    .A1(_3166_),
    .S(_3454_),
    .X(_3457_));
 sky130_fd_sc_hd__clkbuf_1 _7105_ (.A(_3457_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _7106_ (.A0(\mem[8][3] ),
    .A1(_3168_),
    .S(_3454_),
    .X(_3458_));
 sky130_fd_sc_hd__clkbuf_1 _7107_ (.A(_3458_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _7108_ (.A0(\mem[8][4] ),
    .A1(_3170_),
    .S(_3454_),
    .X(_3459_));
 sky130_fd_sc_hd__clkbuf_1 _7109_ (.A(_3459_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _7110_ (.A0(\mem[8][5] ),
    .A1(_3172_),
    .S(_3454_),
    .X(_3460_));
 sky130_fd_sc_hd__clkbuf_1 _7111_ (.A(_3460_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _7112_ (.A0(\mem[8][6] ),
    .A1(_3174_),
    .S(_3454_),
    .X(_3461_));
 sky130_fd_sc_hd__clkbuf_1 _7113_ (.A(_3461_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _7114_ (.A0(\mem[8][7] ),
    .A1(_3176_),
    .S(_3454_),
    .X(_3462_));
 sky130_fd_sc_hd__clkbuf_1 _7115_ (.A(_3462_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _7116_ (.A0(\mem[8][8] ),
    .A1(_3178_),
    .S(_3454_),
    .X(_3463_));
 sky130_fd_sc_hd__clkbuf_1 _7117_ (.A(_3463_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _7118_ (.A0(\mem[8][9] ),
    .A1(_3180_),
    .S(_3454_),
    .X(_3464_));
 sky130_fd_sc_hd__clkbuf_1 _7119_ (.A(_3464_),
    .X(_0265_));
 sky130_fd_sc_hd__buf_6 _7120_ (.A(_3453_),
    .X(_3465_));
 sky130_fd_sc_hd__mux2_1 _7121_ (.A0(\mem[8][10] ),
    .A1(_3182_),
    .S(_3465_),
    .X(_3466_));
 sky130_fd_sc_hd__clkbuf_1 _7122_ (.A(_3466_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _7123_ (.A0(\mem[8][11] ),
    .A1(_3185_),
    .S(_3465_),
    .X(_3467_));
 sky130_fd_sc_hd__clkbuf_1 _7124_ (.A(_3467_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _7125_ (.A0(\mem[8][12] ),
    .A1(_3187_),
    .S(_3465_),
    .X(_3468_));
 sky130_fd_sc_hd__clkbuf_1 _7126_ (.A(_3468_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _7127_ (.A0(\mem[8][13] ),
    .A1(_3189_),
    .S(_3465_),
    .X(_3469_));
 sky130_fd_sc_hd__clkbuf_1 _7128_ (.A(_3469_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _7129_ (.A0(\mem[8][14] ),
    .A1(_3191_),
    .S(_3465_),
    .X(_3470_));
 sky130_fd_sc_hd__clkbuf_1 _7130_ (.A(_3470_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _7131_ (.A0(\mem[8][15] ),
    .A1(_3193_),
    .S(_3465_),
    .X(_3471_));
 sky130_fd_sc_hd__clkbuf_1 _7132_ (.A(_3471_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _7133_ (.A0(\mem[8][16] ),
    .A1(_3195_),
    .S(_3465_),
    .X(_3472_));
 sky130_fd_sc_hd__clkbuf_1 _7134_ (.A(_3472_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _7135_ (.A0(\mem[8][17] ),
    .A1(_3197_),
    .S(_3465_),
    .X(_3473_));
 sky130_fd_sc_hd__clkbuf_1 _7136_ (.A(_3473_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _7137_ (.A0(\mem[8][18] ),
    .A1(_3199_),
    .S(_3465_),
    .X(_3474_));
 sky130_fd_sc_hd__clkbuf_1 _7138_ (.A(_3474_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _7139_ (.A0(\mem[8][19] ),
    .A1(_3201_),
    .S(_3465_),
    .X(_3475_));
 sky130_fd_sc_hd__clkbuf_1 _7140_ (.A(_3475_),
    .X(_0275_));
 sky130_fd_sc_hd__buf_4 _7141_ (.A(_3453_),
    .X(_3476_));
 sky130_fd_sc_hd__mux2_1 _7142_ (.A0(\mem[8][20] ),
    .A1(_3203_),
    .S(_3476_),
    .X(_3477_));
 sky130_fd_sc_hd__clkbuf_1 _7143_ (.A(_3477_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _7144_ (.A0(\mem[8][21] ),
    .A1(_3206_),
    .S(_3476_),
    .X(_3478_));
 sky130_fd_sc_hd__clkbuf_1 _7145_ (.A(_3478_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _7146_ (.A0(\mem[8][22] ),
    .A1(_3208_),
    .S(_3476_),
    .X(_3479_));
 sky130_fd_sc_hd__clkbuf_1 _7147_ (.A(_3479_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _7148_ (.A0(\mem[8][23] ),
    .A1(_3210_),
    .S(_3476_),
    .X(_3480_));
 sky130_fd_sc_hd__clkbuf_1 _7149_ (.A(_3480_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _7150_ (.A0(\mem[8][24] ),
    .A1(_3212_),
    .S(_3476_),
    .X(_3481_));
 sky130_fd_sc_hd__clkbuf_1 _7151_ (.A(_3481_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _7152_ (.A0(\mem[8][25] ),
    .A1(_3214_),
    .S(_3476_),
    .X(_3482_));
 sky130_fd_sc_hd__clkbuf_1 _7153_ (.A(_3482_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _7154_ (.A0(\mem[8][26] ),
    .A1(_3216_),
    .S(_3476_),
    .X(_3483_));
 sky130_fd_sc_hd__clkbuf_1 _7155_ (.A(_3483_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _7156_ (.A0(\mem[8][27] ),
    .A1(_3218_),
    .S(_3476_),
    .X(_3484_));
 sky130_fd_sc_hd__clkbuf_1 _7157_ (.A(_3484_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _7158_ (.A0(\mem[8][28] ),
    .A1(_3220_),
    .S(_3476_),
    .X(_3485_));
 sky130_fd_sc_hd__clkbuf_1 _7159_ (.A(_3485_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _7160_ (.A0(\mem[8][29] ),
    .A1(_3222_),
    .S(_3476_),
    .X(_3486_));
 sky130_fd_sc_hd__clkbuf_1 _7161_ (.A(_3486_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _7162_ (.A0(\mem[8][30] ),
    .A1(_3224_),
    .S(_3453_),
    .X(_3487_));
 sky130_fd_sc_hd__clkbuf_1 _7163_ (.A(_3487_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _7164_ (.A0(\mem[8][31] ),
    .A1(_3226_),
    .S(_3453_),
    .X(_3488_));
 sky130_fd_sc_hd__clkbuf_1 _7165_ (.A(_3488_),
    .X(_0287_));
 sky130_fd_sc_hd__or2b_1 _7166_ (.A(net15),
    .B_N(net16),
    .X(_3489_));
 sky130_fd_sc_hd__or3_4 _7167_ (.A(_3340_),
    .B(_3342_),
    .C(_3489_),
    .X(_3490_));
 sky130_fd_sc_hd__buf_6 _7168_ (.A(_3490_),
    .X(_3491_));
 sky130_fd_sc_hd__mux2_1 _7169_ (.A0(_3086_),
    .A1(\mem[9][0] ),
    .S(_3491_),
    .X(_3492_));
 sky130_fd_sc_hd__clkbuf_1 _7170_ (.A(_3492_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _7171_ (.A0(_3093_),
    .A1(\mem[9][1] ),
    .S(_3491_),
    .X(_3493_));
 sky130_fd_sc_hd__clkbuf_1 _7172_ (.A(_3493_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _7173_ (.A0(_3095_),
    .A1(\mem[9][2] ),
    .S(_3491_),
    .X(_3494_));
 sky130_fd_sc_hd__clkbuf_1 _7174_ (.A(_3494_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _7175_ (.A0(_3097_),
    .A1(\mem[9][3] ),
    .S(_3491_),
    .X(_3495_));
 sky130_fd_sc_hd__clkbuf_1 _7176_ (.A(_3495_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _7177_ (.A0(_3099_),
    .A1(\mem[9][4] ),
    .S(_3491_),
    .X(_3496_));
 sky130_fd_sc_hd__clkbuf_1 _7178_ (.A(_3496_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _7179_ (.A0(_3101_),
    .A1(\mem[9][5] ),
    .S(_3491_),
    .X(_3497_));
 sky130_fd_sc_hd__clkbuf_1 _7180_ (.A(_3497_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _7181_ (.A0(_3103_),
    .A1(\mem[9][6] ),
    .S(_3491_),
    .X(_3498_));
 sky130_fd_sc_hd__clkbuf_1 _7182_ (.A(_3498_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _7183_ (.A0(_3105_),
    .A1(\mem[9][7] ),
    .S(_3491_),
    .X(_3499_));
 sky130_fd_sc_hd__clkbuf_1 _7184_ (.A(_3499_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _7185_ (.A0(_3107_),
    .A1(\mem[9][8] ),
    .S(_3491_),
    .X(_3500_));
 sky130_fd_sc_hd__clkbuf_1 _7186_ (.A(_3500_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _7187_ (.A0(_3109_),
    .A1(\mem[9][9] ),
    .S(_3491_),
    .X(_3501_));
 sky130_fd_sc_hd__clkbuf_1 _7188_ (.A(_3501_),
    .X(_0297_));
 sky130_fd_sc_hd__buf_6 _7189_ (.A(_3490_),
    .X(_3502_));
 sky130_fd_sc_hd__mux2_1 _7190_ (.A0(_3111_),
    .A1(\mem[9][10] ),
    .S(_3502_),
    .X(_3503_));
 sky130_fd_sc_hd__clkbuf_1 _7191_ (.A(_3503_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _7192_ (.A0(_3114_),
    .A1(\mem[9][11] ),
    .S(_3502_),
    .X(_3504_));
 sky130_fd_sc_hd__clkbuf_1 _7193_ (.A(_3504_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _7194_ (.A0(_3116_),
    .A1(\mem[9][12] ),
    .S(_3502_),
    .X(_3505_));
 sky130_fd_sc_hd__clkbuf_1 _7195_ (.A(_3505_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _7196_ (.A0(_3118_),
    .A1(\mem[9][13] ),
    .S(_3502_),
    .X(_3506_));
 sky130_fd_sc_hd__clkbuf_1 _7197_ (.A(_3506_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _7198_ (.A0(_3120_),
    .A1(\mem[9][14] ),
    .S(_3502_),
    .X(_3507_));
 sky130_fd_sc_hd__clkbuf_1 _7199_ (.A(_3507_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _7200_ (.A0(_3122_),
    .A1(\mem[9][15] ),
    .S(_3502_),
    .X(_3508_));
 sky130_fd_sc_hd__clkbuf_1 _7201_ (.A(_3508_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _7202_ (.A0(_3124_),
    .A1(\mem[9][16] ),
    .S(_3502_),
    .X(_3509_));
 sky130_fd_sc_hd__clkbuf_1 _7203_ (.A(_3509_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _7204_ (.A0(_3126_),
    .A1(\mem[9][17] ),
    .S(_3502_),
    .X(_3510_));
 sky130_fd_sc_hd__clkbuf_1 _7205_ (.A(_3510_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _7206_ (.A0(_3128_),
    .A1(\mem[9][18] ),
    .S(_3502_),
    .X(_3511_));
 sky130_fd_sc_hd__clkbuf_1 _7207_ (.A(_3511_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _7208_ (.A0(_3130_),
    .A1(\mem[9][19] ),
    .S(_3502_),
    .X(_3512_));
 sky130_fd_sc_hd__clkbuf_1 _7209_ (.A(_3512_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_4 _7210_ (.A(_3490_),
    .X(_3513_));
 sky130_fd_sc_hd__mux2_1 _7211_ (.A0(_3132_),
    .A1(\mem[9][20] ),
    .S(_3513_),
    .X(_3514_));
 sky130_fd_sc_hd__clkbuf_1 _7212_ (.A(_3514_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _7213_ (.A0(_3135_),
    .A1(\mem[9][21] ),
    .S(_3513_),
    .X(_3515_));
 sky130_fd_sc_hd__clkbuf_1 _7214_ (.A(_3515_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _7215_ (.A0(_3137_),
    .A1(\mem[9][22] ),
    .S(_3513_),
    .X(_3516_));
 sky130_fd_sc_hd__clkbuf_1 _7216_ (.A(_3516_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _7217_ (.A0(_3139_),
    .A1(\mem[9][23] ),
    .S(_3513_),
    .X(_3517_));
 sky130_fd_sc_hd__clkbuf_1 _7218_ (.A(_3517_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _7219_ (.A0(_3141_),
    .A1(\mem[9][24] ),
    .S(_3513_),
    .X(_3518_));
 sky130_fd_sc_hd__clkbuf_1 _7220_ (.A(_3518_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _7221_ (.A0(_3143_),
    .A1(\mem[9][25] ),
    .S(_3513_),
    .X(_3519_));
 sky130_fd_sc_hd__clkbuf_1 _7222_ (.A(_3519_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _7223_ (.A0(_3145_),
    .A1(\mem[9][26] ),
    .S(_3513_),
    .X(_3520_));
 sky130_fd_sc_hd__clkbuf_1 _7224_ (.A(_3520_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _7225_ (.A0(_3147_),
    .A1(\mem[9][27] ),
    .S(_3513_),
    .X(_3521_));
 sky130_fd_sc_hd__clkbuf_1 _7226_ (.A(_3521_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _7227_ (.A0(_3149_),
    .A1(\mem[9][28] ),
    .S(_3513_),
    .X(_3522_));
 sky130_fd_sc_hd__clkbuf_1 _7228_ (.A(_3522_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _7229_ (.A0(_3151_),
    .A1(\mem[9][29] ),
    .S(_3513_),
    .X(_3523_));
 sky130_fd_sc_hd__clkbuf_1 _7230_ (.A(_3523_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _7231_ (.A0(_3153_),
    .A1(\mem[9][30] ),
    .S(_3490_),
    .X(_3524_));
 sky130_fd_sc_hd__clkbuf_1 _7232_ (.A(_3524_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _7233_ (.A0(_3155_),
    .A1(\mem[9][31] ),
    .S(_3490_),
    .X(_3525_));
 sky130_fd_sc_hd__clkbuf_1 _7234_ (.A(_3525_),
    .X(_0319_));
 sky130_fd_sc_hd__or3_4 _7235_ (.A(_3379_),
    .B(_3342_),
    .C(_3489_),
    .X(_3526_));
 sky130_fd_sc_hd__buf_4 _7236_ (.A(_3526_),
    .X(_3527_));
 sky130_fd_sc_hd__mux2_1 _7237_ (.A0(_3086_),
    .A1(\mem[10][0] ),
    .S(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__clkbuf_1 _7238_ (.A(_3528_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _7239_ (.A0(_3093_),
    .A1(\mem[10][1] ),
    .S(_3527_),
    .X(_3529_));
 sky130_fd_sc_hd__clkbuf_1 _7240_ (.A(_3529_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _7241_ (.A0(_3095_),
    .A1(\mem[10][2] ),
    .S(_3527_),
    .X(_3530_));
 sky130_fd_sc_hd__clkbuf_1 _7242_ (.A(_3530_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _7243_ (.A0(_3097_),
    .A1(\mem[10][3] ),
    .S(_3527_),
    .X(_3531_));
 sky130_fd_sc_hd__clkbuf_1 _7244_ (.A(_3531_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _7245_ (.A0(_3099_),
    .A1(\mem[10][4] ),
    .S(_3527_),
    .X(_3532_));
 sky130_fd_sc_hd__clkbuf_1 _7246_ (.A(_3532_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _7247_ (.A0(_3101_),
    .A1(\mem[10][5] ),
    .S(_3527_),
    .X(_3533_));
 sky130_fd_sc_hd__clkbuf_1 _7248_ (.A(_3533_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _7249_ (.A0(_3103_),
    .A1(\mem[10][6] ),
    .S(_3527_),
    .X(_3534_));
 sky130_fd_sc_hd__clkbuf_1 _7250_ (.A(_3534_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _7251_ (.A0(_3105_),
    .A1(\mem[10][7] ),
    .S(_3527_),
    .X(_3535_));
 sky130_fd_sc_hd__clkbuf_1 _7252_ (.A(_3535_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _7253_ (.A0(_3107_),
    .A1(\mem[10][8] ),
    .S(_3527_),
    .X(_3536_));
 sky130_fd_sc_hd__clkbuf_1 _7254_ (.A(_3536_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _7255_ (.A0(_3109_),
    .A1(\mem[10][9] ),
    .S(_3527_),
    .X(_3537_));
 sky130_fd_sc_hd__clkbuf_1 _7256_ (.A(_3537_),
    .X(_0329_));
 sky130_fd_sc_hd__buf_6 _7257_ (.A(_3526_),
    .X(_3538_));
 sky130_fd_sc_hd__mux2_1 _7258_ (.A0(_3111_),
    .A1(\mem[10][10] ),
    .S(_3538_),
    .X(_3539_));
 sky130_fd_sc_hd__clkbuf_1 _7259_ (.A(_3539_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _7260_ (.A0(_3114_),
    .A1(\mem[10][11] ),
    .S(_3538_),
    .X(_3540_));
 sky130_fd_sc_hd__clkbuf_1 _7261_ (.A(_3540_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _7262_ (.A0(_3116_),
    .A1(\mem[10][12] ),
    .S(_3538_),
    .X(_3541_));
 sky130_fd_sc_hd__clkbuf_1 _7263_ (.A(_3541_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _7264_ (.A0(_3118_),
    .A1(\mem[10][13] ),
    .S(_3538_),
    .X(_3542_));
 sky130_fd_sc_hd__clkbuf_1 _7265_ (.A(_3542_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _7266_ (.A0(_3120_),
    .A1(\mem[10][14] ),
    .S(_3538_),
    .X(_3543_));
 sky130_fd_sc_hd__clkbuf_1 _7267_ (.A(_3543_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _7268_ (.A0(_3122_),
    .A1(\mem[10][15] ),
    .S(_3538_),
    .X(_3544_));
 sky130_fd_sc_hd__clkbuf_1 _7269_ (.A(_3544_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _7270_ (.A0(_3124_),
    .A1(\mem[10][16] ),
    .S(_3538_),
    .X(_3545_));
 sky130_fd_sc_hd__clkbuf_1 _7271_ (.A(_3545_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _7272_ (.A0(_3126_),
    .A1(\mem[10][17] ),
    .S(_3538_),
    .X(_3546_));
 sky130_fd_sc_hd__clkbuf_1 _7273_ (.A(_3546_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _7274_ (.A0(_3128_),
    .A1(\mem[10][18] ),
    .S(_3538_),
    .X(_3547_));
 sky130_fd_sc_hd__clkbuf_1 _7275_ (.A(_3547_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _7276_ (.A0(_3130_),
    .A1(\mem[10][19] ),
    .S(_3538_),
    .X(_3548_));
 sky130_fd_sc_hd__clkbuf_1 _7277_ (.A(_3548_),
    .X(_0339_));
 sky130_fd_sc_hd__buf_4 _7278_ (.A(_3526_),
    .X(_3549_));
 sky130_fd_sc_hd__mux2_1 _7279_ (.A0(_3132_),
    .A1(\mem[10][20] ),
    .S(_3549_),
    .X(_3550_));
 sky130_fd_sc_hd__clkbuf_1 _7280_ (.A(_3550_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _7281_ (.A0(_3135_),
    .A1(\mem[10][21] ),
    .S(_3549_),
    .X(_3551_));
 sky130_fd_sc_hd__clkbuf_1 _7282_ (.A(_3551_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _7283_ (.A0(_3137_),
    .A1(\mem[10][22] ),
    .S(_3549_),
    .X(_3552_));
 sky130_fd_sc_hd__clkbuf_1 _7284_ (.A(_3552_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _7285_ (.A0(_3139_),
    .A1(\mem[10][23] ),
    .S(_3549_),
    .X(_3553_));
 sky130_fd_sc_hd__clkbuf_1 _7286_ (.A(_3553_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _7287_ (.A0(_3141_),
    .A1(\mem[10][24] ),
    .S(_3549_),
    .X(_3554_));
 sky130_fd_sc_hd__clkbuf_1 _7288_ (.A(_3554_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _7289_ (.A0(_3143_),
    .A1(\mem[10][25] ),
    .S(_3549_),
    .X(_3555_));
 sky130_fd_sc_hd__clkbuf_1 _7290_ (.A(_3555_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _7291_ (.A0(_3145_),
    .A1(\mem[10][26] ),
    .S(_3549_),
    .X(_3556_));
 sky130_fd_sc_hd__clkbuf_1 _7292_ (.A(_3556_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _7293_ (.A0(_3147_),
    .A1(\mem[10][27] ),
    .S(_3549_),
    .X(_3557_));
 sky130_fd_sc_hd__clkbuf_1 _7294_ (.A(_3557_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _7295_ (.A0(_3149_),
    .A1(\mem[10][28] ),
    .S(_3549_),
    .X(_3558_));
 sky130_fd_sc_hd__clkbuf_1 _7296_ (.A(_3558_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _7297_ (.A0(_3151_),
    .A1(\mem[10][29] ),
    .S(_3549_),
    .X(_3559_));
 sky130_fd_sc_hd__clkbuf_1 _7298_ (.A(_3559_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _7299_ (.A0(_3153_),
    .A1(\mem[10][30] ),
    .S(_3526_),
    .X(_3560_));
 sky130_fd_sc_hd__clkbuf_1 _7300_ (.A(_3560_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _7301_ (.A0(_3155_),
    .A1(\mem[10][31] ),
    .S(_3526_),
    .X(_3561_));
 sky130_fd_sc_hd__clkbuf_1 _7302_ (.A(_3561_),
    .X(_0351_));
 sky130_fd_sc_hd__or3_4 _7303_ (.A(_3088_),
    .B(_3342_),
    .C(_3489_),
    .X(_3562_));
 sky130_fd_sc_hd__buf_6 _7304_ (.A(_3562_),
    .X(_3563_));
 sky130_fd_sc_hd__mux2_1 _7305_ (.A0(_3086_),
    .A1(\mem[11][0] ),
    .S(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__clkbuf_1 _7306_ (.A(_3564_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _7307_ (.A0(_3093_),
    .A1(\mem[11][1] ),
    .S(_3563_),
    .X(_3565_));
 sky130_fd_sc_hd__clkbuf_1 _7308_ (.A(_3565_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _7309_ (.A0(_3095_),
    .A1(\mem[11][2] ),
    .S(_3563_),
    .X(_3566_));
 sky130_fd_sc_hd__clkbuf_1 _7310_ (.A(_3566_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _7311_ (.A0(_3097_),
    .A1(\mem[11][3] ),
    .S(_3563_),
    .X(_3567_));
 sky130_fd_sc_hd__clkbuf_1 _7312_ (.A(_3567_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _7313_ (.A0(_3099_),
    .A1(\mem[11][4] ),
    .S(_3563_),
    .X(_3568_));
 sky130_fd_sc_hd__clkbuf_1 _7314_ (.A(_3568_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _7315_ (.A0(_3101_),
    .A1(\mem[11][5] ),
    .S(_3563_),
    .X(_3569_));
 sky130_fd_sc_hd__clkbuf_1 _7316_ (.A(_3569_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _7317_ (.A0(_3103_),
    .A1(\mem[11][6] ),
    .S(_3563_),
    .X(_3570_));
 sky130_fd_sc_hd__clkbuf_1 _7318_ (.A(_3570_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _7319_ (.A0(_3105_),
    .A1(\mem[11][7] ),
    .S(_3563_),
    .X(_3571_));
 sky130_fd_sc_hd__clkbuf_1 _7320_ (.A(_3571_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _7321_ (.A0(_3107_),
    .A1(\mem[11][8] ),
    .S(_3563_),
    .X(_3572_));
 sky130_fd_sc_hd__clkbuf_1 _7322_ (.A(_3572_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _7323_ (.A0(_3109_),
    .A1(\mem[11][9] ),
    .S(_3563_),
    .X(_3573_));
 sky130_fd_sc_hd__clkbuf_1 _7324_ (.A(_3573_),
    .X(_0361_));
 sky130_fd_sc_hd__buf_6 _7325_ (.A(_3562_),
    .X(_3574_));
 sky130_fd_sc_hd__mux2_1 _7326_ (.A0(_3111_),
    .A1(\mem[11][10] ),
    .S(_3574_),
    .X(_3575_));
 sky130_fd_sc_hd__clkbuf_1 _7327_ (.A(_3575_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _7328_ (.A0(_3114_),
    .A1(\mem[11][11] ),
    .S(_3574_),
    .X(_3576_));
 sky130_fd_sc_hd__clkbuf_1 _7329_ (.A(_3576_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _7330_ (.A0(_3116_),
    .A1(\mem[11][12] ),
    .S(_3574_),
    .X(_3577_));
 sky130_fd_sc_hd__clkbuf_1 _7331_ (.A(_3577_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _7332_ (.A0(_3118_),
    .A1(\mem[11][13] ),
    .S(_3574_),
    .X(_3578_));
 sky130_fd_sc_hd__clkbuf_1 _7333_ (.A(_3578_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _7334_ (.A0(_3120_),
    .A1(\mem[11][14] ),
    .S(_3574_),
    .X(_3579_));
 sky130_fd_sc_hd__clkbuf_1 _7335_ (.A(_3579_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _7336_ (.A0(_3122_),
    .A1(\mem[11][15] ),
    .S(_3574_),
    .X(_3580_));
 sky130_fd_sc_hd__clkbuf_1 _7337_ (.A(_3580_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _7338_ (.A0(_3124_),
    .A1(\mem[11][16] ),
    .S(_3574_),
    .X(_3581_));
 sky130_fd_sc_hd__clkbuf_1 _7339_ (.A(_3581_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _7340_ (.A0(_3126_),
    .A1(\mem[11][17] ),
    .S(_3574_),
    .X(_3582_));
 sky130_fd_sc_hd__clkbuf_1 _7341_ (.A(_3582_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _7342_ (.A0(_3128_),
    .A1(\mem[11][18] ),
    .S(_3574_),
    .X(_3583_));
 sky130_fd_sc_hd__clkbuf_1 _7343_ (.A(_3583_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _7344_ (.A0(_3130_),
    .A1(\mem[11][19] ),
    .S(_3574_),
    .X(_3584_));
 sky130_fd_sc_hd__clkbuf_1 _7345_ (.A(_3584_),
    .X(_0371_));
 sky130_fd_sc_hd__buf_4 _7346_ (.A(_3562_),
    .X(_3585_));
 sky130_fd_sc_hd__mux2_1 _7347_ (.A0(_3132_),
    .A1(\mem[11][20] ),
    .S(_3585_),
    .X(_3586_));
 sky130_fd_sc_hd__clkbuf_1 _7348_ (.A(_3586_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _7349_ (.A0(_3135_),
    .A1(\mem[11][21] ),
    .S(_3585_),
    .X(_3587_));
 sky130_fd_sc_hd__clkbuf_1 _7350_ (.A(_3587_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _7351_ (.A0(_3137_),
    .A1(\mem[11][22] ),
    .S(_3585_),
    .X(_3588_));
 sky130_fd_sc_hd__clkbuf_1 _7352_ (.A(_3588_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _7353_ (.A0(_3139_),
    .A1(\mem[11][23] ),
    .S(_3585_),
    .X(_3589_));
 sky130_fd_sc_hd__clkbuf_1 _7354_ (.A(_3589_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _7355_ (.A0(_3141_),
    .A1(\mem[11][24] ),
    .S(_3585_),
    .X(_3590_));
 sky130_fd_sc_hd__clkbuf_1 _7356_ (.A(_3590_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _7357_ (.A0(_3143_),
    .A1(\mem[11][25] ),
    .S(_3585_),
    .X(_3591_));
 sky130_fd_sc_hd__clkbuf_1 _7358_ (.A(_3591_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _7359_ (.A0(_3145_),
    .A1(\mem[11][26] ),
    .S(_3585_),
    .X(_3592_));
 sky130_fd_sc_hd__clkbuf_1 _7360_ (.A(_3592_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _7361_ (.A0(_3147_),
    .A1(\mem[11][27] ),
    .S(_3585_),
    .X(_3593_));
 sky130_fd_sc_hd__clkbuf_1 _7362_ (.A(_3593_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _7363_ (.A0(_3149_),
    .A1(\mem[11][28] ),
    .S(_3585_),
    .X(_3594_));
 sky130_fd_sc_hd__clkbuf_1 _7364_ (.A(_3594_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _7365_ (.A0(_3151_),
    .A1(\mem[11][29] ),
    .S(_3585_),
    .X(_3595_));
 sky130_fd_sc_hd__clkbuf_1 _7366_ (.A(_3595_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _7367_ (.A0(_3153_),
    .A1(\mem[11][30] ),
    .S(_3562_),
    .X(_3596_));
 sky130_fd_sc_hd__clkbuf_1 _7368_ (.A(_3596_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _7369_ (.A0(_3155_),
    .A1(\mem[11][31] ),
    .S(_3562_),
    .X(_3597_));
 sky130_fd_sc_hd__clkbuf_1 _7370_ (.A(_3597_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _7371_ (.A(net16),
    .B(net15),
    .X(_3598_));
 sky130_fd_sc_hd__and3_2 _7372_ (.A(_3598_),
    .B(_3158_),
    .C(_3302_),
    .X(_3599_));
 sky130_fd_sc_hd__buf_6 _7373_ (.A(_3599_),
    .X(_3600_));
 sky130_fd_sc_hd__mux2_1 _7374_ (.A0(\mem[12][0] ),
    .A1(_3157_),
    .S(_3600_),
    .X(_3601_));
 sky130_fd_sc_hd__clkbuf_1 _7375_ (.A(_3601_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _7376_ (.A0(\mem[12][1] ),
    .A1(_3164_),
    .S(_3600_),
    .X(_3602_));
 sky130_fd_sc_hd__clkbuf_1 _7377_ (.A(_3602_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _7378_ (.A0(\mem[12][2] ),
    .A1(_3166_),
    .S(_3600_),
    .X(_3603_));
 sky130_fd_sc_hd__clkbuf_1 _7379_ (.A(_3603_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _7380_ (.A0(\mem[12][3] ),
    .A1(_3168_),
    .S(_3600_),
    .X(_3604_));
 sky130_fd_sc_hd__clkbuf_1 _7381_ (.A(_3604_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _7382_ (.A0(\mem[12][4] ),
    .A1(_3170_),
    .S(_3600_),
    .X(_3605_));
 sky130_fd_sc_hd__clkbuf_1 _7383_ (.A(_3605_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _7384_ (.A0(\mem[12][5] ),
    .A1(_3172_),
    .S(_3600_),
    .X(_3606_));
 sky130_fd_sc_hd__clkbuf_1 _7385_ (.A(_3606_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _7386_ (.A0(\mem[12][6] ),
    .A1(_3174_),
    .S(_3600_),
    .X(_3607_));
 sky130_fd_sc_hd__clkbuf_1 _7387_ (.A(_3607_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _7388_ (.A0(\mem[12][7] ),
    .A1(_3176_),
    .S(_3600_),
    .X(_3608_));
 sky130_fd_sc_hd__clkbuf_1 _7389_ (.A(_3608_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _7390_ (.A0(\mem[12][8] ),
    .A1(_3178_),
    .S(_3600_),
    .X(_3609_));
 sky130_fd_sc_hd__clkbuf_1 _7391_ (.A(_3609_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _7392_ (.A0(\mem[12][9] ),
    .A1(_3180_),
    .S(_3600_),
    .X(_3610_));
 sky130_fd_sc_hd__clkbuf_1 _7393_ (.A(_3610_),
    .X(_0393_));
 sky130_fd_sc_hd__buf_6 _7394_ (.A(_3599_),
    .X(_3611_));
 sky130_fd_sc_hd__mux2_1 _7395_ (.A0(\mem[12][10] ),
    .A1(_3182_),
    .S(_3611_),
    .X(_3612_));
 sky130_fd_sc_hd__clkbuf_1 _7396_ (.A(_3612_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _7397_ (.A0(\mem[12][11] ),
    .A1(_3185_),
    .S(_3611_),
    .X(_3613_));
 sky130_fd_sc_hd__clkbuf_1 _7398_ (.A(_3613_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _7399_ (.A0(\mem[12][12] ),
    .A1(_3187_),
    .S(_3611_),
    .X(_3614_));
 sky130_fd_sc_hd__clkbuf_1 _7400_ (.A(_3614_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _7401_ (.A0(\mem[12][13] ),
    .A1(_3189_),
    .S(_3611_),
    .X(_3615_));
 sky130_fd_sc_hd__clkbuf_1 _7402_ (.A(_3615_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _7403_ (.A0(\mem[12][14] ),
    .A1(_3191_),
    .S(_3611_),
    .X(_3616_));
 sky130_fd_sc_hd__clkbuf_1 _7404_ (.A(_3616_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _7405_ (.A0(\mem[12][15] ),
    .A1(_3193_),
    .S(_3611_),
    .X(_3617_));
 sky130_fd_sc_hd__clkbuf_1 _7406_ (.A(_3617_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _7407_ (.A0(\mem[12][16] ),
    .A1(_3195_),
    .S(_3611_),
    .X(_3618_));
 sky130_fd_sc_hd__clkbuf_1 _7408_ (.A(_3618_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _7409_ (.A0(\mem[12][17] ),
    .A1(_3197_),
    .S(_3611_),
    .X(_3619_));
 sky130_fd_sc_hd__clkbuf_1 _7410_ (.A(_3619_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _7411_ (.A0(\mem[12][18] ),
    .A1(_3199_),
    .S(_3611_),
    .X(_3620_));
 sky130_fd_sc_hd__clkbuf_1 _7412_ (.A(_3620_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _7413_ (.A0(\mem[12][19] ),
    .A1(_3201_),
    .S(_3611_),
    .X(_3621_));
 sky130_fd_sc_hd__clkbuf_1 _7414_ (.A(_3621_),
    .X(_0403_));
 sky130_fd_sc_hd__buf_4 _7415_ (.A(_3599_),
    .X(_3622_));
 sky130_fd_sc_hd__mux2_1 _7416_ (.A0(\mem[12][20] ),
    .A1(_3203_),
    .S(_3622_),
    .X(_3623_));
 sky130_fd_sc_hd__clkbuf_1 _7417_ (.A(_3623_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _7418_ (.A0(\mem[12][21] ),
    .A1(_3206_),
    .S(_3622_),
    .X(_3624_));
 sky130_fd_sc_hd__clkbuf_1 _7419_ (.A(_3624_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _7420_ (.A0(\mem[12][22] ),
    .A1(_3208_),
    .S(_3622_),
    .X(_3625_));
 sky130_fd_sc_hd__clkbuf_1 _7421_ (.A(_3625_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _7422_ (.A0(\mem[12][23] ),
    .A1(_3210_),
    .S(_3622_),
    .X(_3626_));
 sky130_fd_sc_hd__clkbuf_1 _7423_ (.A(_3626_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _7424_ (.A0(\mem[12][24] ),
    .A1(_3212_),
    .S(_3622_),
    .X(_3627_));
 sky130_fd_sc_hd__clkbuf_1 _7425_ (.A(_3627_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _7426_ (.A0(\mem[12][25] ),
    .A1(_3214_),
    .S(_3622_),
    .X(_3628_));
 sky130_fd_sc_hd__clkbuf_1 _7427_ (.A(_3628_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _7428_ (.A0(\mem[12][26] ),
    .A1(_3216_),
    .S(_3622_),
    .X(_3629_));
 sky130_fd_sc_hd__clkbuf_1 _7429_ (.A(_3629_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _7430_ (.A0(\mem[12][27] ),
    .A1(_3218_),
    .S(_3622_),
    .X(_3630_));
 sky130_fd_sc_hd__clkbuf_1 _7431_ (.A(_3630_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _7432_ (.A0(\mem[12][28] ),
    .A1(_3220_),
    .S(_3622_),
    .X(_3631_));
 sky130_fd_sc_hd__clkbuf_1 _7433_ (.A(_3631_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _7434_ (.A0(\mem[12][29] ),
    .A1(_3222_),
    .S(_3622_),
    .X(_3632_));
 sky130_fd_sc_hd__clkbuf_1 _7435_ (.A(_3632_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _7436_ (.A0(\mem[12][30] ),
    .A1(_3224_),
    .S(_3599_),
    .X(_3633_));
 sky130_fd_sc_hd__clkbuf_1 _7437_ (.A(_3633_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _7438_ (.A0(\mem[12][31] ),
    .A1(_3226_),
    .S(_3599_),
    .X(_3634_));
 sky130_fd_sc_hd__clkbuf_1 _7439_ (.A(_3634_),
    .X(_0415_));
 sky130_fd_sc_hd__and4_2 _7440_ (.A(net16),
    .B(net15),
    .C(_3158_),
    .D(_3159_),
    .X(_3635_));
 sky130_fd_sc_hd__buf_4 _7441_ (.A(_3635_),
    .X(_3636_));
 sky130_fd_sc_hd__mux2_1 _7442_ (.A0(\mem[13][0] ),
    .A1(_3157_),
    .S(_3636_),
    .X(_3637_));
 sky130_fd_sc_hd__clkbuf_1 _7443_ (.A(_3637_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _7444_ (.A0(\mem[13][1] ),
    .A1(_3164_),
    .S(_3636_),
    .X(_3638_));
 sky130_fd_sc_hd__clkbuf_1 _7445_ (.A(_3638_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _7446_ (.A0(\mem[13][2] ),
    .A1(_3166_),
    .S(_3636_),
    .X(_3639_));
 sky130_fd_sc_hd__clkbuf_1 _7447_ (.A(_3639_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _7448_ (.A0(\mem[13][3] ),
    .A1(_3168_),
    .S(_3636_),
    .X(_3640_));
 sky130_fd_sc_hd__clkbuf_1 _7449_ (.A(_3640_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _7450_ (.A0(\mem[13][4] ),
    .A1(_3170_),
    .S(_3636_),
    .X(_3641_));
 sky130_fd_sc_hd__clkbuf_1 _7451_ (.A(_3641_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _7452_ (.A0(\mem[13][5] ),
    .A1(_3172_),
    .S(_3636_),
    .X(_3642_));
 sky130_fd_sc_hd__clkbuf_1 _7453_ (.A(_3642_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _7454_ (.A0(\mem[13][6] ),
    .A1(_3174_),
    .S(_3636_),
    .X(_3643_));
 sky130_fd_sc_hd__clkbuf_1 _7455_ (.A(_3643_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _7456_ (.A0(\mem[13][7] ),
    .A1(_3176_),
    .S(_3636_),
    .X(_3644_));
 sky130_fd_sc_hd__clkbuf_1 _7457_ (.A(_3644_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _7458_ (.A0(\mem[13][8] ),
    .A1(_3178_),
    .S(_3636_),
    .X(_3645_));
 sky130_fd_sc_hd__clkbuf_1 _7459_ (.A(_3645_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _7460_ (.A0(\mem[13][9] ),
    .A1(_3180_),
    .S(_3636_),
    .X(_3646_));
 sky130_fd_sc_hd__clkbuf_1 _7461_ (.A(_3646_),
    .X(_0425_));
 sky130_fd_sc_hd__buf_4 _7462_ (.A(_3635_),
    .X(_3647_));
 sky130_fd_sc_hd__mux2_1 _7463_ (.A0(\mem[13][10] ),
    .A1(_3182_),
    .S(_3647_),
    .X(_3648_));
 sky130_fd_sc_hd__clkbuf_1 _7464_ (.A(_3648_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _7465_ (.A0(\mem[13][11] ),
    .A1(_3185_),
    .S(_3647_),
    .X(_3649_));
 sky130_fd_sc_hd__clkbuf_1 _7466_ (.A(_3649_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _7467_ (.A0(\mem[13][12] ),
    .A1(_3187_),
    .S(_3647_),
    .X(_3650_));
 sky130_fd_sc_hd__clkbuf_1 _7468_ (.A(_3650_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _7469_ (.A0(\mem[13][13] ),
    .A1(_3189_),
    .S(_3647_),
    .X(_3651_));
 sky130_fd_sc_hd__clkbuf_1 _7470_ (.A(_3651_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _7471_ (.A0(\mem[13][14] ),
    .A1(_3191_),
    .S(_3647_),
    .X(_3652_));
 sky130_fd_sc_hd__clkbuf_1 _7472_ (.A(_3652_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _7473_ (.A0(\mem[13][15] ),
    .A1(_3193_),
    .S(_3647_),
    .X(_3653_));
 sky130_fd_sc_hd__clkbuf_1 _7474_ (.A(_3653_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _7475_ (.A0(\mem[13][16] ),
    .A1(_3195_),
    .S(_3647_),
    .X(_3654_));
 sky130_fd_sc_hd__clkbuf_1 _7476_ (.A(_3654_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _7477_ (.A0(\mem[13][17] ),
    .A1(_3197_),
    .S(_3647_),
    .X(_3655_));
 sky130_fd_sc_hd__clkbuf_1 _7478_ (.A(_3655_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _7479_ (.A0(\mem[13][18] ),
    .A1(_3199_),
    .S(_3647_),
    .X(_3656_));
 sky130_fd_sc_hd__clkbuf_1 _7480_ (.A(_3656_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _7481_ (.A0(\mem[13][19] ),
    .A1(_3201_),
    .S(_3647_),
    .X(_3657_));
 sky130_fd_sc_hd__clkbuf_1 _7482_ (.A(_3657_),
    .X(_0435_));
 sky130_fd_sc_hd__buf_4 _7483_ (.A(_3635_),
    .X(_3658_));
 sky130_fd_sc_hd__mux2_1 _7484_ (.A0(\mem[13][20] ),
    .A1(_3203_),
    .S(_3658_),
    .X(_3659_));
 sky130_fd_sc_hd__clkbuf_1 _7485_ (.A(_3659_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _7486_ (.A0(\mem[13][21] ),
    .A1(_3206_),
    .S(_3658_),
    .X(_3660_));
 sky130_fd_sc_hd__clkbuf_1 _7487_ (.A(_3660_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _7488_ (.A0(\mem[13][22] ),
    .A1(_3208_),
    .S(_3658_),
    .X(_3661_));
 sky130_fd_sc_hd__clkbuf_1 _7489_ (.A(_3661_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _7490_ (.A0(\mem[13][23] ),
    .A1(_3210_),
    .S(_3658_),
    .X(_3662_));
 sky130_fd_sc_hd__clkbuf_1 _7491_ (.A(_3662_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _7492_ (.A0(\mem[13][24] ),
    .A1(_3212_),
    .S(_3658_),
    .X(_3663_));
 sky130_fd_sc_hd__clkbuf_1 _7493_ (.A(_3663_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _7494_ (.A0(\mem[13][25] ),
    .A1(_3214_),
    .S(_3658_),
    .X(_3664_));
 sky130_fd_sc_hd__clkbuf_1 _7495_ (.A(_3664_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _7496_ (.A0(\mem[13][26] ),
    .A1(_3216_),
    .S(_3658_),
    .X(_3665_));
 sky130_fd_sc_hd__clkbuf_1 _7497_ (.A(_3665_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _7498_ (.A0(\mem[13][27] ),
    .A1(_3218_),
    .S(_3658_),
    .X(_3666_));
 sky130_fd_sc_hd__clkbuf_1 _7499_ (.A(_3666_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _7500_ (.A0(\mem[13][28] ),
    .A1(_3220_),
    .S(_3658_),
    .X(_3667_));
 sky130_fd_sc_hd__clkbuf_1 _7501_ (.A(_3667_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _7502_ (.A0(\mem[13][29] ),
    .A1(_3222_),
    .S(_3658_),
    .X(_3668_));
 sky130_fd_sc_hd__clkbuf_1 _7503_ (.A(_3668_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _7504_ (.A0(\mem[13][30] ),
    .A1(_3224_),
    .S(_3635_),
    .X(_3669_));
 sky130_fd_sc_hd__clkbuf_1 _7505_ (.A(_3669_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _7506_ (.A0(\mem[13][31] ),
    .A1(_3226_),
    .S(_3635_),
    .X(_3670_));
 sky130_fd_sc_hd__clkbuf_1 _7507_ (.A(_3670_),
    .X(_0447_));
 sky130_fd_sc_hd__or3_4 _7508_ (.A(_3089_),
    .B(_3379_),
    .C(_3342_),
    .X(_3671_));
 sky130_fd_sc_hd__buf_6 _7509_ (.A(_3671_),
    .X(_3672_));
 sky130_fd_sc_hd__mux2_1 _7510_ (.A0(_3086_),
    .A1(\mem[14][0] ),
    .S(_3672_),
    .X(_3673_));
 sky130_fd_sc_hd__clkbuf_1 _7511_ (.A(_3673_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _7512_ (.A0(_3093_),
    .A1(\mem[14][1] ),
    .S(_3672_),
    .X(_3674_));
 sky130_fd_sc_hd__clkbuf_1 _7513_ (.A(_3674_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _7514_ (.A0(_3095_),
    .A1(\mem[14][2] ),
    .S(_3672_),
    .X(_3675_));
 sky130_fd_sc_hd__clkbuf_1 _7515_ (.A(_3675_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _7516_ (.A0(_3097_),
    .A1(\mem[14][3] ),
    .S(_3672_),
    .X(_3676_));
 sky130_fd_sc_hd__clkbuf_1 _7517_ (.A(_3676_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _7518_ (.A0(_3099_),
    .A1(\mem[14][4] ),
    .S(_3672_),
    .X(_3677_));
 sky130_fd_sc_hd__clkbuf_1 _7519_ (.A(_3677_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _7520_ (.A0(_3101_),
    .A1(\mem[14][5] ),
    .S(_3672_),
    .X(_3678_));
 sky130_fd_sc_hd__clkbuf_1 _7521_ (.A(_3678_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _7522_ (.A0(_3103_),
    .A1(\mem[14][6] ),
    .S(_3672_),
    .X(_3679_));
 sky130_fd_sc_hd__clkbuf_1 _7523_ (.A(_3679_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _7524_ (.A0(_3105_),
    .A1(\mem[14][7] ),
    .S(_3672_),
    .X(_3680_));
 sky130_fd_sc_hd__clkbuf_1 _7525_ (.A(_3680_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _7526_ (.A0(_3107_),
    .A1(\mem[14][8] ),
    .S(_3672_),
    .X(_3681_));
 sky130_fd_sc_hd__clkbuf_1 _7527_ (.A(_3681_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _7528_ (.A0(_3109_),
    .A1(\mem[14][9] ),
    .S(_3672_),
    .X(_3682_));
 sky130_fd_sc_hd__clkbuf_1 _7529_ (.A(_3682_),
    .X(_0457_));
 sky130_fd_sc_hd__buf_6 _7530_ (.A(_3671_),
    .X(_3683_));
 sky130_fd_sc_hd__mux2_1 _7531_ (.A0(_3111_),
    .A1(\mem[14][10] ),
    .S(_3683_),
    .X(_3684_));
 sky130_fd_sc_hd__clkbuf_1 _7532_ (.A(_3684_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _7533_ (.A0(_3114_),
    .A1(\mem[14][11] ),
    .S(_3683_),
    .X(_3685_));
 sky130_fd_sc_hd__clkbuf_1 _7534_ (.A(_3685_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _7535_ (.A0(_3116_),
    .A1(\mem[14][12] ),
    .S(_3683_),
    .X(_3686_));
 sky130_fd_sc_hd__clkbuf_1 _7536_ (.A(_3686_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _7537_ (.A0(_3118_),
    .A1(\mem[14][13] ),
    .S(_3683_),
    .X(_3687_));
 sky130_fd_sc_hd__clkbuf_1 _7538_ (.A(_3687_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _7539_ (.A0(_3120_),
    .A1(\mem[14][14] ),
    .S(_3683_),
    .X(_3688_));
 sky130_fd_sc_hd__clkbuf_1 _7540_ (.A(_3688_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _7541_ (.A0(_3122_),
    .A1(\mem[14][15] ),
    .S(_3683_),
    .X(_3689_));
 sky130_fd_sc_hd__clkbuf_1 _7542_ (.A(_3689_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _7543_ (.A0(_3124_),
    .A1(\mem[14][16] ),
    .S(_3683_),
    .X(_3690_));
 sky130_fd_sc_hd__clkbuf_1 _7544_ (.A(_3690_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _7545_ (.A0(_3126_),
    .A1(\mem[14][17] ),
    .S(_3683_),
    .X(_3691_));
 sky130_fd_sc_hd__clkbuf_1 _7546_ (.A(_3691_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _7547_ (.A0(_3128_),
    .A1(\mem[14][18] ),
    .S(_3683_),
    .X(_3692_));
 sky130_fd_sc_hd__clkbuf_1 _7548_ (.A(_3692_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _7549_ (.A0(_3130_),
    .A1(\mem[14][19] ),
    .S(_3683_),
    .X(_3693_));
 sky130_fd_sc_hd__clkbuf_1 _7550_ (.A(_3693_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_4 _7551_ (.A(_3671_),
    .X(_3694_));
 sky130_fd_sc_hd__mux2_1 _7552_ (.A0(_3132_),
    .A1(\mem[14][20] ),
    .S(_3694_),
    .X(_3695_));
 sky130_fd_sc_hd__clkbuf_1 _7553_ (.A(_3695_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _7554_ (.A0(_3135_),
    .A1(\mem[14][21] ),
    .S(_3694_),
    .X(_3696_));
 sky130_fd_sc_hd__clkbuf_1 _7555_ (.A(_3696_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _7556_ (.A0(_3137_),
    .A1(\mem[14][22] ),
    .S(_3694_),
    .X(_3697_));
 sky130_fd_sc_hd__clkbuf_1 _7557_ (.A(_3697_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _7558_ (.A0(_3139_),
    .A1(\mem[14][23] ),
    .S(_3694_),
    .X(_3698_));
 sky130_fd_sc_hd__clkbuf_1 _7559_ (.A(_3698_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _7560_ (.A0(_3141_),
    .A1(\mem[14][24] ),
    .S(_3694_),
    .X(_3699_));
 sky130_fd_sc_hd__clkbuf_1 _7561_ (.A(_3699_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _7562_ (.A0(_3143_),
    .A1(\mem[14][25] ),
    .S(_3694_),
    .X(_3700_));
 sky130_fd_sc_hd__clkbuf_1 _7563_ (.A(_3700_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _7564_ (.A0(_3145_),
    .A1(\mem[14][26] ),
    .S(_3694_),
    .X(_3701_));
 sky130_fd_sc_hd__clkbuf_1 _7565_ (.A(_3701_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _7566_ (.A0(_3147_),
    .A1(\mem[14][27] ),
    .S(_3694_),
    .X(_3702_));
 sky130_fd_sc_hd__clkbuf_1 _7567_ (.A(_3702_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _7568_ (.A0(_3149_),
    .A1(\mem[14][28] ),
    .S(_3694_),
    .X(_3703_));
 sky130_fd_sc_hd__clkbuf_1 _7569_ (.A(_3703_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _7570_ (.A0(_3151_),
    .A1(\mem[14][29] ),
    .S(_3694_),
    .X(_3704_));
 sky130_fd_sc_hd__clkbuf_1 _7571_ (.A(_3704_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _7572_ (.A0(_3153_),
    .A1(\mem[14][30] ),
    .S(_3671_),
    .X(_3705_));
 sky130_fd_sc_hd__clkbuf_1 _7573_ (.A(_3705_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _7574_ (.A0(_3155_),
    .A1(\mem[14][31] ),
    .S(_3671_),
    .X(_3706_));
 sky130_fd_sc_hd__clkbuf_1 _7575_ (.A(_3706_),
    .X(_0479_));
 sky130_fd_sc_hd__and4_2 _7576_ (.A(net14),
    .B(net13),
    .C(_3598_),
    .D(_3158_),
    .X(_3707_));
 sky130_fd_sc_hd__buf_4 _7577_ (.A(_3707_),
    .X(_3708_));
 sky130_fd_sc_hd__mux2_1 _7578_ (.A0(\mem[15][0] ),
    .A1(_3157_),
    .S(_3708_),
    .X(_3709_));
 sky130_fd_sc_hd__clkbuf_1 _7579_ (.A(_3709_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _7580_ (.A0(\mem[15][1] ),
    .A1(_3164_),
    .S(_3708_),
    .X(_3710_));
 sky130_fd_sc_hd__clkbuf_1 _7581_ (.A(_3710_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _7582_ (.A0(\mem[15][2] ),
    .A1(_3166_),
    .S(_3708_),
    .X(_3711_));
 sky130_fd_sc_hd__clkbuf_1 _7583_ (.A(_3711_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _7584_ (.A0(\mem[15][3] ),
    .A1(_3168_),
    .S(_3708_),
    .X(_3712_));
 sky130_fd_sc_hd__clkbuf_1 _7585_ (.A(_3712_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _7586_ (.A0(\mem[15][4] ),
    .A1(_3170_),
    .S(_3708_),
    .X(_3713_));
 sky130_fd_sc_hd__clkbuf_1 _7587_ (.A(_3713_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _7588_ (.A0(\mem[15][5] ),
    .A1(_3172_),
    .S(_3708_),
    .X(_3714_));
 sky130_fd_sc_hd__clkbuf_1 _7589_ (.A(_3714_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _7590_ (.A0(\mem[15][6] ),
    .A1(_3174_),
    .S(_3708_),
    .X(_3715_));
 sky130_fd_sc_hd__clkbuf_1 _7591_ (.A(_3715_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _7592_ (.A0(\mem[15][7] ),
    .A1(_3176_),
    .S(_3708_),
    .X(_3716_));
 sky130_fd_sc_hd__clkbuf_1 _7593_ (.A(_3716_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _7594_ (.A0(\mem[15][8] ),
    .A1(_3178_),
    .S(_3708_),
    .X(_3717_));
 sky130_fd_sc_hd__clkbuf_1 _7595_ (.A(_3717_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _7596_ (.A0(\mem[15][9] ),
    .A1(_3180_),
    .S(_3708_),
    .X(_3718_));
 sky130_fd_sc_hd__clkbuf_1 _7597_ (.A(_3718_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_4 _7598_ (.A(_3707_),
    .X(_3719_));
 sky130_fd_sc_hd__mux2_1 _7599_ (.A0(\mem[15][10] ),
    .A1(_3182_),
    .S(_3719_),
    .X(_3720_));
 sky130_fd_sc_hd__clkbuf_1 _7600_ (.A(_3720_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _7601_ (.A0(\mem[15][11] ),
    .A1(_3185_),
    .S(_3719_),
    .X(_3721_));
 sky130_fd_sc_hd__clkbuf_1 _7602_ (.A(_3721_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _7603_ (.A0(\mem[15][12] ),
    .A1(_3187_),
    .S(_3719_),
    .X(_3722_));
 sky130_fd_sc_hd__clkbuf_1 _7604_ (.A(_3722_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _7605_ (.A0(\mem[15][13] ),
    .A1(_3189_),
    .S(_3719_),
    .X(_3723_));
 sky130_fd_sc_hd__clkbuf_1 _7606_ (.A(_3723_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _7607_ (.A0(\mem[15][14] ),
    .A1(_3191_),
    .S(_3719_),
    .X(_3724_));
 sky130_fd_sc_hd__clkbuf_1 _7608_ (.A(_3724_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _7609_ (.A0(\mem[15][15] ),
    .A1(_3193_),
    .S(_3719_),
    .X(_3725_));
 sky130_fd_sc_hd__clkbuf_1 _7610_ (.A(_3725_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _7611_ (.A0(\mem[15][16] ),
    .A1(_3195_),
    .S(_3719_),
    .X(_3726_));
 sky130_fd_sc_hd__clkbuf_1 _7612_ (.A(_3726_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _7613_ (.A0(\mem[15][17] ),
    .A1(_3197_),
    .S(_3719_),
    .X(_3727_));
 sky130_fd_sc_hd__clkbuf_1 _7614_ (.A(_3727_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _7615_ (.A0(\mem[15][18] ),
    .A1(_3199_),
    .S(_3719_),
    .X(_3728_));
 sky130_fd_sc_hd__clkbuf_1 _7616_ (.A(_3728_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _7617_ (.A0(\mem[15][19] ),
    .A1(_3201_),
    .S(_3719_),
    .X(_3729_));
 sky130_fd_sc_hd__clkbuf_1 _7618_ (.A(_3729_),
    .X(_0499_));
 sky130_fd_sc_hd__buf_4 _7619_ (.A(_3707_),
    .X(_3730_));
 sky130_fd_sc_hd__mux2_1 _7620_ (.A0(\mem[15][20] ),
    .A1(_3203_),
    .S(_3730_),
    .X(_3731_));
 sky130_fd_sc_hd__clkbuf_1 _7621_ (.A(_3731_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _7622_ (.A0(\mem[15][21] ),
    .A1(_3206_),
    .S(_3730_),
    .X(_3732_));
 sky130_fd_sc_hd__clkbuf_1 _7623_ (.A(_3732_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _7624_ (.A0(\mem[15][22] ),
    .A1(_3208_),
    .S(_3730_),
    .X(_3733_));
 sky130_fd_sc_hd__clkbuf_1 _7625_ (.A(_3733_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _7626_ (.A0(\mem[15][23] ),
    .A1(_3210_),
    .S(_3730_),
    .X(_3734_));
 sky130_fd_sc_hd__clkbuf_1 _7627_ (.A(_3734_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _7628_ (.A0(\mem[15][24] ),
    .A1(_3212_),
    .S(_3730_),
    .X(_3735_));
 sky130_fd_sc_hd__clkbuf_1 _7629_ (.A(_3735_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _7630_ (.A0(\mem[15][25] ),
    .A1(_3214_),
    .S(_3730_),
    .X(_3736_));
 sky130_fd_sc_hd__clkbuf_1 _7631_ (.A(_3736_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _7632_ (.A0(\mem[15][26] ),
    .A1(_3216_),
    .S(_3730_),
    .X(_3737_));
 sky130_fd_sc_hd__clkbuf_1 _7633_ (.A(_3737_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _7634_ (.A0(\mem[15][27] ),
    .A1(_3218_),
    .S(_3730_),
    .X(_3738_));
 sky130_fd_sc_hd__clkbuf_1 _7635_ (.A(_3738_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _7636_ (.A0(\mem[15][28] ),
    .A1(_3220_),
    .S(_3730_),
    .X(_3739_));
 sky130_fd_sc_hd__clkbuf_1 _7637_ (.A(_3739_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _7638_ (.A0(\mem[15][29] ),
    .A1(_3222_),
    .S(_3730_),
    .X(_3740_));
 sky130_fd_sc_hd__clkbuf_1 _7639_ (.A(_3740_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _7640_ (.A0(\mem[15][30] ),
    .A1(_3224_),
    .S(_3707_),
    .X(_3741_));
 sky130_fd_sc_hd__clkbuf_1 _7641_ (.A(_3741_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _7642_ (.A0(\mem[15][31] ),
    .A1(_3226_),
    .S(_3707_),
    .X(_3742_));
 sky130_fd_sc_hd__clkbuf_1 _7643_ (.A(_3742_),
    .X(_0511_));
 sky130_fd_sc_hd__buf_2 _7644_ (.A(net18),
    .X(_3743_));
 sky130_fd_sc_hd__and2_1 _7645_ (.A(net17),
    .B(net12),
    .X(_3744_));
 sky130_fd_sc_hd__clkbuf_2 _7646_ (.A(_3744_),
    .X(_3745_));
 sky130_fd_sc_hd__and3_4 _7647_ (.A(_3745_),
    .B(_3160_),
    .C(_3302_),
    .X(_3746_));
 sky130_fd_sc_hd__buf_6 _7648_ (.A(_3746_),
    .X(_3747_));
 sky130_fd_sc_hd__mux2_1 _7649_ (.A0(\mem[16][0] ),
    .A1(_3743_),
    .S(_3747_),
    .X(_3748_));
 sky130_fd_sc_hd__clkbuf_1 _7650_ (.A(_3748_),
    .X(_0512_));
 sky130_fd_sc_hd__buf_2 _7651_ (.A(net29),
    .X(_3749_));
 sky130_fd_sc_hd__mux2_1 _7652_ (.A0(\mem[16][1] ),
    .A1(_3749_),
    .S(_3747_),
    .X(_3750_));
 sky130_fd_sc_hd__clkbuf_1 _7653_ (.A(_3750_),
    .X(_0513_));
 sky130_fd_sc_hd__buf_2 _7654_ (.A(net40),
    .X(_3751_));
 sky130_fd_sc_hd__mux2_1 _7655_ (.A0(\mem[16][2] ),
    .A1(_3751_),
    .S(_3747_),
    .X(_3752_));
 sky130_fd_sc_hd__clkbuf_1 _7656_ (.A(_3752_),
    .X(_0514_));
 sky130_fd_sc_hd__buf_2 _7657_ (.A(net43),
    .X(_3753_));
 sky130_fd_sc_hd__mux2_1 _7658_ (.A0(\mem[16][3] ),
    .A1(_3753_),
    .S(_3747_),
    .X(_3754_));
 sky130_fd_sc_hd__clkbuf_1 _7659_ (.A(_3754_),
    .X(_0515_));
 sky130_fd_sc_hd__buf_2 _7660_ (.A(net44),
    .X(_3755_));
 sky130_fd_sc_hd__mux2_1 _7661_ (.A0(\mem[16][4] ),
    .A1(_3755_),
    .S(_3747_),
    .X(_3756_));
 sky130_fd_sc_hd__clkbuf_1 _7662_ (.A(_3756_),
    .X(_0516_));
 sky130_fd_sc_hd__buf_2 _7663_ (.A(net45),
    .X(_3757_));
 sky130_fd_sc_hd__mux2_1 _7664_ (.A0(\mem[16][5] ),
    .A1(_3757_),
    .S(_3747_),
    .X(_3758_));
 sky130_fd_sc_hd__clkbuf_1 _7665_ (.A(_3758_),
    .X(_0517_));
 sky130_fd_sc_hd__buf_2 _7666_ (.A(net46),
    .X(_3759_));
 sky130_fd_sc_hd__mux2_1 _7667_ (.A0(\mem[16][6] ),
    .A1(_3759_),
    .S(_3747_),
    .X(_3760_));
 sky130_fd_sc_hd__clkbuf_1 _7668_ (.A(_3760_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_2 _7669_ (.A(net47),
    .X(_3761_));
 sky130_fd_sc_hd__mux2_1 _7670_ (.A0(\mem[16][7] ),
    .A1(_3761_),
    .S(_3747_),
    .X(_3762_));
 sky130_fd_sc_hd__clkbuf_1 _7671_ (.A(_3762_),
    .X(_0519_));
 sky130_fd_sc_hd__buf_2 _7672_ (.A(net48),
    .X(_3763_));
 sky130_fd_sc_hd__mux2_1 _7673_ (.A0(\mem[16][8] ),
    .A1(_3763_),
    .S(_3747_),
    .X(_3764_));
 sky130_fd_sc_hd__clkbuf_1 _7674_ (.A(_3764_),
    .X(_0520_));
 sky130_fd_sc_hd__buf_2 _7675_ (.A(net49),
    .X(_3765_));
 sky130_fd_sc_hd__mux2_1 _7676_ (.A0(\mem[16][9] ),
    .A1(_3765_),
    .S(_3747_),
    .X(_3766_));
 sky130_fd_sc_hd__clkbuf_1 _7677_ (.A(_3766_),
    .X(_0521_));
 sky130_fd_sc_hd__buf_2 _7678_ (.A(net19),
    .X(_3767_));
 sky130_fd_sc_hd__buf_6 _7679_ (.A(_3746_),
    .X(_3768_));
 sky130_fd_sc_hd__mux2_1 _7680_ (.A0(\mem[16][10] ),
    .A1(_3767_),
    .S(_3768_),
    .X(_3769_));
 sky130_fd_sc_hd__clkbuf_1 _7681_ (.A(_3769_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_2 _7682_ (.A(net20),
    .X(_3770_));
 sky130_fd_sc_hd__mux2_1 _7683_ (.A0(\mem[16][11] ),
    .A1(_3770_),
    .S(_3768_),
    .X(_3771_));
 sky130_fd_sc_hd__clkbuf_1 _7684_ (.A(_3771_),
    .X(_0523_));
 sky130_fd_sc_hd__buf_2 _7685_ (.A(net21),
    .X(_3772_));
 sky130_fd_sc_hd__mux2_1 _7686_ (.A0(\mem[16][12] ),
    .A1(_3772_),
    .S(_3768_),
    .X(_3773_));
 sky130_fd_sc_hd__clkbuf_1 _7687_ (.A(_3773_),
    .X(_0524_));
 sky130_fd_sc_hd__buf_2 _7688_ (.A(net22),
    .X(_3774_));
 sky130_fd_sc_hd__mux2_1 _7689_ (.A0(\mem[16][13] ),
    .A1(_3774_),
    .S(_3768_),
    .X(_3775_));
 sky130_fd_sc_hd__clkbuf_1 _7690_ (.A(_3775_),
    .X(_0525_));
 sky130_fd_sc_hd__buf_2 _7691_ (.A(net23),
    .X(_3776_));
 sky130_fd_sc_hd__mux2_1 _7692_ (.A0(\mem[16][14] ),
    .A1(_3776_),
    .S(_3768_),
    .X(_3777_));
 sky130_fd_sc_hd__clkbuf_1 _7693_ (.A(_3777_),
    .X(_0526_));
 sky130_fd_sc_hd__buf_2 _7694_ (.A(net24),
    .X(_3778_));
 sky130_fd_sc_hd__mux2_1 _7695_ (.A0(\mem[16][15] ),
    .A1(_3778_),
    .S(_3768_),
    .X(_3779_));
 sky130_fd_sc_hd__clkbuf_1 _7696_ (.A(_3779_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _7697_ (.A(net25),
    .X(_3780_));
 sky130_fd_sc_hd__mux2_1 _7698_ (.A0(\mem[16][16] ),
    .A1(_3780_),
    .S(_3768_),
    .X(_3781_));
 sky130_fd_sc_hd__clkbuf_1 _7699_ (.A(_3781_),
    .X(_0528_));
 sky130_fd_sc_hd__buf_2 _7700_ (.A(net26),
    .X(_3782_));
 sky130_fd_sc_hd__mux2_1 _7701_ (.A0(\mem[16][17] ),
    .A1(_3782_),
    .S(_3768_),
    .X(_3783_));
 sky130_fd_sc_hd__clkbuf_1 _7702_ (.A(_3783_),
    .X(_0529_));
 sky130_fd_sc_hd__buf_2 _7703_ (.A(net27),
    .X(_3784_));
 sky130_fd_sc_hd__mux2_1 _7704_ (.A0(\mem[16][18] ),
    .A1(_3784_),
    .S(_3768_),
    .X(_3785_));
 sky130_fd_sc_hd__clkbuf_1 _7705_ (.A(_3785_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_2 _7706_ (.A(net28),
    .X(_3786_));
 sky130_fd_sc_hd__mux2_1 _7707_ (.A0(\mem[16][19] ),
    .A1(_3786_),
    .S(_3768_),
    .X(_3787_));
 sky130_fd_sc_hd__clkbuf_1 _7708_ (.A(_3787_),
    .X(_0531_));
 sky130_fd_sc_hd__buf_2 _7709_ (.A(net30),
    .X(_3788_));
 sky130_fd_sc_hd__buf_4 _7710_ (.A(_3746_),
    .X(_3789_));
 sky130_fd_sc_hd__mux2_1 _7711_ (.A0(\mem[16][20] ),
    .A1(_3788_),
    .S(_3789_),
    .X(_3790_));
 sky130_fd_sc_hd__clkbuf_1 _7712_ (.A(_3790_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_4 _7713_ (.A(net31),
    .X(_3791_));
 sky130_fd_sc_hd__mux2_1 _7714_ (.A0(\mem[16][21] ),
    .A1(_3791_),
    .S(_3789_),
    .X(_3792_));
 sky130_fd_sc_hd__clkbuf_1 _7715_ (.A(_3792_),
    .X(_0533_));
 sky130_fd_sc_hd__buf_2 _7716_ (.A(net32),
    .X(_3793_));
 sky130_fd_sc_hd__mux2_1 _7717_ (.A0(\mem[16][22] ),
    .A1(_3793_),
    .S(_3789_),
    .X(_3794_));
 sky130_fd_sc_hd__clkbuf_1 _7718_ (.A(_3794_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_4 _7719_ (.A(net33),
    .X(_3795_));
 sky130_fd_sc_hd__mux2_1 _7720_ (.A0(\mem[16][23] ),
    .A1(_3795_),
    .S(_3789_),
    .X(_3796_));
 sky130_fd_sc_hd__clkbuf_1 _7721_ (.A(_3796_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _7722_ (.A(net34),
    .X(_3797_));
 sky130_fd_sc_hd__mux2_1 _7723_ (.A0(\mem[16][24] ),
    .A1(_3797_),
    .S(_3789_),
    .X(_3798_));
 sky130_fd_sc_hd__clkbuf_1 _7724_ (.A(_3798_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_2 _7725_ (.A(net35),
    .X(_3799_));
 sky130_fd_sc_hd__mux2_1 _7726_ (.A0(\mem[16][25] ),
    .A1(_3799_),
    .S(_3789_),
    .X(_3800_));
 sky130_fd_sc_hd__clkbuf_1 _7727_ (.A(_3800_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_2 _7728_ (.A(net36),
    .X(_3801_));
 sky130_fd_sc_hd__mux2_1 _7729_ (.A0(\mem[16][26] ),
    .A1(_3801_),
    .S(_3789_),
    .X(_3802_));
 sky130_fd_sc_hd__clkbuf_1 _7730_ (.A(_3802_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_2 _7731_ (.A(net37),
    .X(_3803_));
 sky130_fd_sc_hd__mux2_1 _7732_ (.A0(\mem[16][27] ),
    .A1(_3803_),
    .S(_3789_),
    .X(_3804_));
 sky130_fd_sc_hd__clkbuf_1 _7733_ (.A(_3804_),
    .X(_0539_));
 sky130_fd_sc_hd__buf_2 _7734_ (.A(net38),
    .X(_3805_));
 sky130_fd_sc_hd__mux2_1 _7735_ (.A0(\mem[16][28] ),
    .A1(_3805_),
    .S(_3789_),
    .X(_3806_));
 sky130_fd_sc_hd__clkbuf_1 _7736_ (.A(_3806_),
    .X(_0540_));
 sky130_fd_sc_hd__buf_2 _7737_ (.A(net39),
    .X(_3807_));
 sky130_fd_sc_hd__mux2_1 _7738_ (.A0(\mem[16][29] ),
    .A1(_3807_),
    .S(_3789_),
    .X(_3808_));
 sky130_fd_sc_hd__clkbuf_1 _7739_ (.A(_3808_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_4 _7740_ (.A(net41),
    .X(_3809_));
 sky130_fd_sc_hd__mux2_1 _7741_ (.A0(\mem[16][30] ),
    .A1(_3809_),
    .S(_3746_),
    .X(_3810_));
 sky130_fd_sc_hd__clkbuf_1 _7742_ (.A(_3810_),
    .X(_0542_));
 sky130_fd_sc_hd__buf_2 _7743_ (.A(net42),
    .X(_3811_));
 sky130_fd_sc_hd__mux2_1 _7744_ (.A0(\mem[16][31] ),
    .A1(_3811_),
    .S(_3746_),
    .X(_3812_));
 sky130_fd_sc_hd__clkbuf_1 _7745_ (.A(_3812_),
    .X(_0543_));
 sky130_fd_sc_hd__and3_4 _7746_ (.A(_3745_),
    .B(_3159_),
    .C(_3160_),
    .X(_3813_));
 sky130_fd_sc_hd__buf_6 _7747_ (.A(_3813_),
    .X(_3814_));
 sky130_fd_sc_hd__mux2_1 _7748_ (.A0(\mem[17][0] ),
    .A1(_3743_),
    .S(_3814_),
    .X(_3815_));
 sky130_fd_sc_hd__clkbuf_1 _7749_ (.A(_3815_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _7750_ (.A0(\mem[17][1] ),
    .A1(_3749_),
    .S(_3814_),
    .X(_3816_));
 sky130_fd_sc_hd__clkbuf_1 _7751_ (.A(_3816_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _7752_ (.A0(\mem[17][2] ),
    .A1(_3751_),
    .S(_3814_),
    .X(_3817_));
 sky130_fd_sc_hd__clkbuf_1 _7753_ (.A(_3817_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _7754_ (.A0(\mem[17][3] ),
    .A1(_3753_),
    .S(_3814_),
    .X(_3818_));
 sky130_fd_sc_hd__clkbuf_1 _7755_ (.A(_3818_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _7756_ (.A0(\mem[17][4] ),
    .A1(_3755_),
    .S(_3814_),
    .X(_3819_));
 sky130_fd_sc_hd__clkbuf_1 _7757_ (.A(_3819_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _7758_ (.A0(\mem[17][5] ),
    .A1(_3757_),
    .S(_3814_),
    .X(_3820_));
 sky130_fd_sc_hd__clkbuf_1 _7759_ (.A(_3820_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _7760_ (.A0(\mem[17][6] ),
    .A1(_3759_),
    .S(_3814_),
    .X(_3821_));
 sky130_fd_sc_hd__clkbuf_1 _7761_ (.A(_3821_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _7762_ (.A0(\mem[17][7] ),
    .A1(_3761_),
    .S(_3814_),
    .X(_3822_));
 sky130_fd_sc_hd__clkbuf_1 _7763_ (.A(_3822_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _7764_ (.A0(\mem[17][8] ),
    .A1(_3763_),
    .S(_3814_),
    .X(_3823_));
 sky130_fd_sc_hd__clkbuf_1 _7765_ (.A(_3823_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _7766_ (.A0(\mem[17][9] ),
    .A1(_3765_),
    .S(_3814_),
    .X(_3824_));
 sky130_fd_sc_hd__clkbuf_1 _7767_ (.A(_3824_),
    .X(_0553_));
 sky130_fd_sc_hd__buf_6 _7768_ (.A(_3813_),
    .X(_3825_));
 sky130_fd_sc_hd__mux2_1 _7769_ (.A0(\mem[17][10] ),
    .A1(_3767_),
    .S(_3825_),
    .X(_3826_));
 sky130_fd_sc_hd__clkbuf_1 _7770_ (.A(_3826_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _7771_ (.A0(\mem[17][11] ),
    .A1(_3770_),
    .S(_3825_),
    .X(_3827_));
 sky130_fd_sc_hd__clkbuf_1 _7772_ (.A(_3827_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _7773_ (.A0(\mem[17][12] ),
    .A1(_3772_),
    .S(_3825_),
    .X(_3828_));
 sky130_fd_sc_hd__clkbuf_1 _7774_ (.A(_3828_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _7775_ (.A0(\mem[17][13] ),
    .A1(_3774_),
    .S(_3825_),
    .X(_3829_));
 sky130_fd_sc_hd__clkbuf_1 _7776_ (.A(_3829_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _7777_ (.A0(\mem[17][14] ),
    .A1(_3776_),
    .S(_3825_),
    .X(_3830_));
 sky130_fd_sc_hd__clkbuf_1 _7778_ (.A(_3830_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _7779_ (.A0(\mem[17][15] ),
    .A1(_3778_),
    .S(_3825_),
    .X(_3831_));
 sky130_fd_sc_hd__clkbuf_1 _7780_ (.A(_3831_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _7781_ (.A0(\mem[17][16] ),
    .A1(_3780_),
    .S(_3825_),
    .X(_3832_));
 sky130_fd_sc_hd__clkbuf_1 _7782_ (.A(_3832_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _7783_ (.A0(\mem[17][17] ),
    .A1(_3782_),
    .S(_3825_),
    .X(_3833_));
 sky130_fd_sc_hd__clkbuf_1 _7784_ (.A(_3833_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _7785_ (.A0(\mem[17][18] ),
    .A1(_3784_),
    .S(_3825_),
    .X(_3834_));
 sky130_fd_sc_hd__clkbuf_1 _7786_ (.A(_3834_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _7787_ (.A0(\mem[17][19] ),
    .A1(_3786_),
    .S(_3825_),
    .X(_3835_));
 sky130_fd_sc_hd__clkbuf_1 _7788_ (.A(_3835_),
    .X(_0563_));
 sky130_fd_sc_hd__buf_4 _7789_ (.A(_3813_),
    .X(_3836_));
 sky130_fd_sc_hd__mux2_1 _7790_ (.A0(\mem[17][20] ),
    .A1(_3788_),
    .S(_3836_),
    .X(_3837_));
 sky130_fd_sc_hd__clkbuf_1 _7791_ (.A(_3837_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _7792_ (.A0(\mem[17][21] ),
    .A1(_3791_),
    .S(_3836_),
    .X(_3838_));
 sky130_fd_sc_hd__clkbuf_1 _7793_ (.A(_3838_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _7794_ (.A0(\mem[17][22] ),
    .A1(_3793_),
    .S(_3836_),
    .X(_3839_));
 sky130_fd_sc_hd__clkbuf_1 _7795_ (.A(_3839_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _7796_ (.A0(\mem[17][23] ),
    .A1(_3795_),
    .S(_3836_),
    .X(_3840_));
 sky130_fd_sc_hd__clkbuf_1 _7797_ (.A(_3840_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _7798_ (.A0(\mem[17][24] ),
    .A1(_3797_),
    .S(_3836_),
    .X(_3841_));
 sky130_fd_sc_hd__clkbuf_1 _7799_ (.A(_3841_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _7800_ (.A0(\mem[17][25] ),
    .A1(_3799_),
    .S(_3836_),
    .X(_3842_));
 sky130_fd_sc_hd__clkbuf_1 _7801_ (.A(_3842_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _7802_ (.A0(\mem[17][26] ),
    .A1(_3801_),
    .S(_3836_),
    .X(_3843_));
 sky130_fd_sc_hd__clkbuf_1 _7803_ (.A(_3843_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _7804_ (.A0(\mem[17][27] ),
    .A1(_3803_),
    .S(_3836_),
    .X(_3844_));
 sky130_fd_sc_hd__clkbuf_1 _7805_ (.A(_3844_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _7806_ (.A0(\mem[17][28] ),
    .A1(_3805_),
    .S(_3836_),
    .X(_3845_));
 sky130_fd_sc_hd__clkbuf_1 _7807_ (.A(_3845_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _7808_ (.A0(\mem[17][29] ),
    .A1(_3807_),
    .S(_3836_),
    .X(_3846_));
 sky130_fd_sc_hd__clkbuf_1 _7809_ (.A(_3846_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _7810_ (.A0(\mem[17][30] ),
    .A1(_3809_),
    .S(_3813_),
    .X(_3847_));
 sky130_fd_sc_hd__clkbuf_1 _7811_ (.A(_3847_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _7812_ (.A0(\mem[17][31] ),
    .A1(_3811_),
    .S(_3813_),
    .X(_3848_));
 sky130_fd_sc_hd__clkbuf_1 _7813_ (.A(_3848_),
    .X(_0575_));
 sky130_fd_sc_hd__and3_2 _7814_ (.A(_3745_),
    .B(_3160_),
    .C(_3228_),
    .X(_3849_));
 sky130_fd_sc_hd__buf_4 _7815_ (.A(_3849_),
    .X(_3850_));
 sky130_fd_sc_hd__mux2_1 _7816_ (.A0(\mem[18][0] ),
    .A1(_3743_),
    .S(_3850_),
    .X(_3851_));
 sky130_fd_sc_hd__clkbuf_1 _7817_ (.A(_3851_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _7818_ (.A0(\mem[18][1] ),
    .A1(_3749_),
    .S(_3850_),
    .X(_3852_));
 sky130_fd_sc_hd__clkbuf_1 _7819_ (.A(_3852_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _7820_ (.A0(\mem[18][2] ),
    .A1(_3751_),
    .S(_3850_),
    .X(_3853_));
 sky130_fd_sc_hd__clkbuf_1 _7821_ (.A(_3853_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _7822_ (.A0(\mem[18][3] ),
    .A1(_3753_),
    .S(_3850_),
    .X(_3854_));
 sky130_fd_sc_hd__clkbuf_1 _7823_ (.A(_3854_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _7824_ (.A0(\mem[18][4] ),
    .A1(_3755_),
    .S(_3850_),
    .X(_3855_));
 sky130_fd_sc_hd__clkbuf_1 _7825_ (.A(_3855_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _7826_ (.A0(\mem[18][5] ),
    .A1(_3757_),
    .S(_3850_),
    .X(_3856_));
 sky130_fd_sc_hd__clkbuf_1 _7827_ (.A(_3856_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _7828_ (.A0(\mem[18][6] ),
    .A1(_3759_),
    .S(_3850_),
    .X(_3857_));
 sky130_fd_sc_hd__clkbuf_1 _7829_ (.A(_3857_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _7830_ (.A0(\mem[18][7] ),
    .A1(_3761_),
    .S(_3850_),
    .X(_3858_));
 sky130_fd_sc_hd__clkbuf_1 _7831_ (.A(_3858_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _7832_ (.A0(\mem[18][8] ),
    .A1(_3763_),
    .S(_3850_),
    .X(_3859_));
 sky130_fd_sc_hd__clkbuf_1 _7833_ (.A(_3859_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _7834_ (.A0(\mem[18][9] ),
    .A1(_3765_),
    .S(_3850_),
    .X(_3860_));
 sky130_fd_sc_hd__clkbuf_1 _7835_ (.A(_3860_),
    .X(_0585_));
 sky130_fd_sc_hd__buf_6 _7836_ (.A(_3849_),
    .X(_3861_));
 sky130_fd_sc_hd__mux2_1 _7837_ (.A0(\mem[18][10] ),
    .A1(_3767_),
    .S(_3861_),
    .X(_3862_));
 sky130_fd_sc_hd__clkbuf_1 _7838_ (.A(_3862_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _7839_ (.A0(\mem[18][11] ),
    .A1(_3770_),
    .S(_3861_),
    .X(_3863_));
 sky130_fd_sc_hd__clkbuf_1 _7840_ (.A(_3863_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _7841_ (.A0(\mem[18][12] ),
    .A1(_3772_),
    .S(_3861_),
    .X(_3864_));
 sky130_fd_sc_hd__clkbuf_1 _7842_ (.A(_3864_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _7843_ (.A0(\mem[18][13] ),
    .A1(_3774_),
    .S(_3861_),
    .X(_3865_));
 sky130_fd_sc_hd__clkbuf_1 _7844_ (.A(_3865_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _7845_ (.A0(\mem[18][14] ),
    .A1(_3776_),
    .S(_3861_),
    .X(_3866_));
 sky130_fd_sc_hd__clkbuf_1 _7846_ (.A(_3866_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _7847_ (.A0(\mem[18][15] ),
    .A1(_3778_),
    .S(_3861_),
    .X(_3867_));
 sky130_fd_sc_hd__clkbuf_1 _7848_ (.A(_3867_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _7849_ (.A0(\mem[18][16] ),
    .A1(_3780_),
    .S(_3861_),
    .X(_3868_));
 sky130_fd_sc_hd__clkbuf_1 _7850_ (.A(_3868_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _7851_ (.A0(\mem[18][17] ),
    .A1(_3782_),
    .S(_3861_),
    .X(_3869_));
 sky130_fd_sc_hd__clkbuf_1 _7852_ (.A(_3869_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _7853_ (.A0(\mem[18][18] ),
    .A1(_3784_),
    .S(_3861_),
    .X(_3870_));
 sky130_fd_sc_hd__clkbuf_1 _7854_ (.A(_3870_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _7855_ (.A0(\mem[18][19] ),
    .A1(_3786_),
    .S(_3861_),
    .X(_3871_));
 sky130_fd_sc_hd__clkbuf_1 _7856_ (.A(_3871_),
    .X(_0595_));
 sky130_fd_sc_hd__buf_4 _7857_ (.A(_3849_),
    .X(_3872_));
 sky130_fd_sc_hd__mux2_1 _7858_ (.A0(\mem[18][20] ),
    .A1(_3788_),
    .S(_3872_),
    .X(_3873_));
 sky130_fd_sc_hd__clkbuf_1 _7859_ (.A(_3873_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _7860_ (.A0(\mem[18][21] ),
    .A1(_3791_),
    .S(_3872_),
    .X(_3874_));
 sky130_fd_sc_hd__clkbuf_1 _7861_ (.A(_3874_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _7862_ (.A0(\mem[18][22] ),
    .A1(_3793_),
    .S(_3872_),
    .X(_3875_));
 sky130_fd_sc_hd__clkbuf_1 _7863_ (.A(_3875_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _7864_ (.A0(\mem[18][23] ),
    .A1(_3795_),
    .S(_3872_),
    .X(_3876_));
 sky130_fd_sc_hd__clkbuf_1 _7865_ (.A(_3876_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _7866_ (.A0(\mem[18][24] ),
    .A1(_3797_),
    .S(_3872_),
    .X(_3877_));
 sky130_fd_sc_hd__clkbuf_1 _7867_ (.A(_3877_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _7868_ (.A0(\mem[18][25] ),
    .A1(_3799_),
    .S(_3872_),
    .X(_3878_));
 sky130_fd_sc_hd__clkbuf_1 _7869_ (.A(_3878_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _7870_ (.A0(\mem[18][26] ),
    .A1(_3801_),
    .S(_3872_),
    .X(_3879_));
 sky130_fd_sc_hd__clkbuf_1 _7871_ (.A(_3879_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _7872_ (.A0(\mem[18][27] ),
    .A1(_3803_),
    .S(_3872_),
    .X(_3880_));
 sky130_fd_sc_hd__clkbuf_1 _7873_ (.A(_3880_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _7874_ (.A0(\mem[18][28] ),
    .A1(_3805_),
    .S(_3872_),
    .X(_3881_));
 sky130_fd_sc_hd__clkbuf_1 _7875_ (.A(_3881_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _7876_ (.A0(\mem[18][29] ),
    .A1(_3807_),
    .S(_3872_),
    .X(_3882_));
 sky130_fd_sc_hd__clkbuf_1 _7877_ (.A(_3882_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _7878_ (.A0(\mem[18][30] ),
    .A1(_3809_),
    .S(_3849_),
    .X(_3883_));
 sky130_fd_sc_hd__clkbuf_1 _7879_ (.A(_3883_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _7880_ (.A0(\mem[18][31] ),
    .A1(_3811_),
    .S(_3849_),
    .X(_3884_));
 sky130_fd_sc_hd__clkbuf_1 _7881_ (.A(_3884_),
    .X(_0607_));
 sky130_fd_sc_hd__and4_4 _7882_ (.A(net14),
    .B(net13),
    .C(_3744_),
    .D(_3160_),
    .X(_3885_));
 sky130_fd_sc_hd__buf_6 _7883_ (.A(_3885_),
    .X(_3886_));
 sky130_fd_sc_hd__mux2_1 _7884_ (.A0(\mem[19][0] ),
    .A1(_3743_),
    .S(_3886_),
    .X(_3887_));
 sky130_fd_sc_hd__clkbuf_1 _7885_ (.A(_3887_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _7886_ (.A0(\mem[19][1] ),
    .A1(_3749_),
    .S(_3886_),
    .X(_3888_));
 sky130_fd_sc_hd__clkbuf_1 _7887_ (.A(_3888_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _7888_ (.A0(\mem[19][2] ),
    .A1(_3751_),
    .S(_3886_),
    .X(_3889_));
 sky130_fd_sc_hd__clkbuf_1 _7889_ (.A(_3889_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _7890_ (.A0(\mem[19][3] ),
    .A1(_3753_),
    .S(_3886_),
    .X(_3890_));
 sky130_fd_sc_hd__clkbuf_1 _7891_ (.A(_3890_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _7892_ (.A0(\mem[19][4] ),
    .A1(_3755_),
    .S(_3886_),
    .X(_3891_));
 sky130_fd_sc_hd__clkbuf_1 _7893_ (.A(_3891_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _7894_ (.A0(\mem[19][5] ),
    .A1(_3757_),
    .S(_3886_),
    .X(_3892_));
 sky130_fd_sc_hd__clkbuf_1 _7895_ (.A(_3892_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _7896_ (.A0(\mem[19][6] ),
    .A1(_3759_),
    .S(_3886_),
    .X(_3893_));
 sky130_fd_sc_hd__clkbuf_1 _7897_ (.A(_3893_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _7898_ (.A0(\mem[19][7] ),
    .A1(_3761_),
    .S(_3886_),
    .X(_3894_));
 sky130_fd_sc_hd__clkbuf_1 _7899_ (.A(_3894_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _7900_ (.A0(\mem[19][8] ),
    .A1(_3763_),
    .S(_3886_),
    .X(_3895_));
 sky130_fd_sc_hd__clkbuf_1 _7901_ (.A(_3895_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _7902_ (.A0(\mem[19][9] ),
    .A1(_3765_),
    .S(_3886_),
    .X(_3896_));
 sky130_fd_sc_hd__clkbuf_1 _7903_ (.A(_3896_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_6 _7904_ (.A(_3885_),
    .X(_3897_));
 sky130_fd_sc_hd__mux2_1 _7905_ (.A0(\mem[19][10] ),
    .A1(_3767_),
    .S(_3897_),
    .X(_3898_));
 sky130_fd_sc_hd__clkbuf_1 _7906_ (.A(_3898_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _7907_ (.A0(\mem[19][11] ),
    .A1(_3770_),
    .S(_3897_),
    .X(_3899_));
 sky130_fd_sc_hd__clkbuf_1 _7908_ (.A(_3899_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _7909_ (.A0(\mem[19][12] ),
    .A1(_3772_),
    .S(_3897_),
    .X(_3900_));
 sky130_fd_sc_hd__clkbuf_1 _7910_ (.A(_3900_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _7911_ (.A0(\mem[19][13] ),
    .A1(_3774_),
    .S(_3897_),
    .X(_3901_));
 sky130_fd_sc_hd__clkbuf_1 _7912_ (.A(_3901_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _7913_ (.A0(\mem[19][14] ),
    .A1(_3776_),
    .S(_3897_),
    .X(_3902_));
 sky130_fd_sc_hd__clkbuf_1 _7914_ (.A(_3902_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _7915_ (.A0(\mem[19][15] ),
    .A1(_3778_),
    .S(_3897_),
    .X(_3903_));
 sky130_fd_sc_hd__clkbuf_1 _7916_ (.A(_3903_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _7917_ (.A0(\mem[19][16] ),
    .A1(_3780_),
    .S(_3897_),
    .X(_3904_));
 sky130_fd_sc_hd__clkbuf_1 _7918_ (.A(_3904_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _7919_ (.A0(\mem[19][17] ),
    .A1(_3782_),
    .S(_3897_),
    .X(_3905_));
 sky130_fd_sc_hd__clkbuf_1 _7920_ (.A(_3905_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _7921_ (.A0(\mem[19][18] ),
    .A1(_3784_),
    .S(_3897_),
    .X(_3906_));
 sky130_fd_sc_hd__clkbuf_1 _7922_ (.A(_3906_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _7923_ (.A0(\mem[19][19] ),
    .A1(_3786_),
    .S(_3897_),
    .X(_3907_));
 sky130_fd_sc_hd__clkbuf_1 _7924_ (.A(_3907_),
    .X(_0627_));
 sky130_fd_sc_hd__buf_4 _7925_ (.A(_3885_),
    .X(_3908_));
 sky130_fd_sc_hd__mux2_1 _7926_ (.A0(\mem[19][20] ),
    .A1(_3788_),
    .S(_3908_),
    .X(_3909_));
 sky130_fd_sc_hd__clkbuf_1 _7927_ (.A(_3909_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _7928_ (.A0(\mem[19][21] ),
    .A1(_3791_),
    .S(_3908_),
    .X(_3910_));
 sky130_fd_sc_hd__clkbuf_1 _7929_ (.A(_3910_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _7930_ (.A0(\mem[19][22] ),
    .A1(_3793_),
    .S(_3908_),
    .X(_3911_));
 sky130_fd_sc_hd__clkbuf_1 _7931_ (.A(_3911_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _7932_ (.A0(\mem[19][23] ),
    .A1(_3795_),
    .S(_3908_),
    .X(_3912_));
 sky130_fd_sc_hd__clkbuf_1 _7933_ (.A(_3912_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _7934_ (.A0(\mem[19][24] ),
    .A1(_3797_),
    .S(_3908_),
    .X(_3913_));
 sky130_fd_sc_hd__clkbuf_1 _7935_ (.A(_3913_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _7936_ (.A0(\mem[19][25] ),
    .A1(_3799_),
    .S(_3908_),
    .X(_3914_));
 sky130_fd_sc_hd__clkbuf_1 _7937_ (.A(_3914_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _7938_ (.A0(\mem[19][26] ),
    .A1(_3801_),
    .S(_3908_),
    .X(_3915_));
 sky130_fd_sc_hd__clkbuf_1 _7939_ (.A(_3915_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _7940_ (.A0(\mem[19][27] ),
    .A1(_3803_),
    .S(_3908_),
    .X(_3916_));
 sky130_fd_sc_hd__clkbuf_1 _7941_ (.A(_3916_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _7942_ (.A0(\mem[19][28] ),
    .A1(_3805_),
    .S(_3908_),
    .X(_3917_));
 sky130_fd_sc_hd__clkbuf_1 _7943_ (.A(_3917_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _7944_ (.A0(\mem[19][29] ),
    .A1(_3807_),
    .S(_3908_),
    .X(_3918_));
 sky130_fd_sc_hd__clkbuf_1 _7945_ (.A(_3918_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _7946_ (.A0(\mem[19][30] ),
    .A1(_3809_),
    .S(_3885_),
    .X(_3919_));
 sky130_fd_sc_hd__clkbuf_1 _7947_ (.A(_3919_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _7948_ (.A0(\mem[19][31] ),
    .A1(_3811_),
    .S(_3885_),
    .X(_3920_));
 sky130_fd_sc_hd__clkbuf_1 _7949_ (.A(_3920_),
    .X(_0639_));
 sky130_fd_sc_hd__and3_2 _7950_ (.A(_3745_),
    .B(_3302_),
    .C(_3303_),
    .X(_3921_));
 sky130_fd_sc_hd__clkbuf_8 _7951_ (.A(_3921_),
    .X(_3922_));
 sky130_fd_sc_hd__mux2_1 _7952_ (.A0(\mem[20][0] ),
    .A1(_3743_),
    .S(_3922_),
    .X(_3923_));
 sky130_fd_sc_hd__clkbuf_1 _7953_ (.A(_3923_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _7954_ (.A0(\mem[20][1] ),
    .A1(_3749_),
    .S(_3922_),
    .X(_3924_));
 sky130_fd_sc_hd__clkbuf_1 _7955_ (.A(_3924_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _7956_ (.A0(\mem[20][2] ),
    .A1(_3751_),
    .S(_3922_),
    .X(_3925_));
 sky130_fd_sc_hd__clkbuf_1 _7957_ (.A(_3925_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _7958_ (.A0(\mem[20][3] ),
    .A1(_3753_),
    .S(_3922_),
    .X(_3926_));
 sky130_fd_sc_hd__clkbuf_1 _7959_ (.A(_3926_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _7960_ (.A0(\mem[20][4] ),
    .A1(_3755_),
    .S(_3922_),
    .X(_3927_));
 sky130_fd_sc_hd__clkbuf_1 _7961_ (.A(_3927_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _7962_ (.A0(\mem[20][5] ),
    .A1(_3757_),
    .S(_3922_),
    .X(_3928_));
 sky130_fd_sc_hd__clkbuf_1 _7963_ (.A(_3928_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _7964_ (.A0(\mem[20][6] ),
    .A1(_3759_),
    .S(_3922_),
    .X(_3929_));
 sky130_fd_sc_hd__clkbuf_1 _7965_ (.A(_3929_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _7966_ (.A0(\mem[20][7] ),
    .A1(_3761_),
    .S(_3922_),
    .X(_3930_));
 sky130_fd_sc_hd__clkbuf_1 _7967_ (.A(_3930_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _7968_ (.A0(\mem[20][8] ),
    .A1(_3763_),
    .S(_3922_),
    .X(_3931_));
 sky130_fd_sc_hd__clkbuf_1 _7969_ (.A(_3931_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _7970_ (.A0(\mem[20][9] ),
    .A1(_3765_),
    .S(_3922_),
    .X(_3932_));
 sky130_fd_sc_hd__clkbuf_1 _7971_ (.A(_3932_),
    .X(_0649_));
 sky130_fd_sc_hd__buf_6 _7972_ (.A(_3921_),
    .X(_3933_));
 sky130_fd_sc_hd__mux2_1 _7973_ (.A0(\mem[20][10] ),
    .A1(_3767_),
    .S(_3933_),
    .X(_3934_));
 sky130_fd_sc_hd__clkbuf_1 _7974_ (.A(_3934_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _7975_ (.A0(\mem[20][11] ),
    .A1(_3770_),
    .S(_3933_),
    .X(_3935_));
 sky130_fd_sc_hd__clkbuf_1 _7976_ (.A(_3935_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _7977_ (.A0(\mem[20][12] ),
    .A1(_3772_),
    .S(_3933_),
    .X(_3936_));
 sky130_fd_sc_hd__clkbuf_1 _7978_ (.A(_3936_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _7979_ (.A0(\mem[20][13] ),
    .A1(_3774_),
    .S(_3933_),
    .X(_3937_));
 sky130_fd_sc_hd__clkbuf_1 _7980_ (.A(_3937_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _7981_ (.A0(\mem[20][14] ),
    .A1(_3776_),
    .S(_3933_),
    .X(_3938_));
 sky130_fd_sc_hd__clkbuf_1 _7982_ (.A(_3938_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _7983_ (.A0(\mem[20][15] ),
    .A1(_3778_),
    .S(_3933_),
    .X(_3939_));
 sky130_fd_sc_hd__clkbuf_1 _7984_ (.A(_3939_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _7985_ (.A0(\mem[20][16] ),
    .A1(_3780_),
    .S(_3933_),
    .X(_3940_));
 sky130_fd_sc_hd__clkbuf_1 _7986_ (.A(_3940_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _7987_ (.A0(\mem[20][17] ),
    .A1(_3782_),
    .S(_3933_),
    .X(_3941_));
 sky130_fd_sc_hd__clkbuf_1 _7988_ (.A(_3941_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _7989_ (.A0(\mem[20][18] ),
    .A1(_3784_),
    .S(_3933_),
    .X(_3942_));
 sky130_fd_sc_hd__clkbuf_1 _7990_ (.A(_3942_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _7991_ (.A0(\mem[20][19] ),
    .A1(_3786_),
    .S(_3933_),
    .X(_3943_));
 sky130_fd_sc_hd__clkbuf_1 _7992_ (.A(_3943_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_4 _7993_ (.A(_3921_),
    .X(_3944_));
 sky130_fd_sc_hd__mux2_1 _7994_ (.A0(\mem[20][20] ),
    .A1(_3788_),
    .S(_3944_),
    .X(_3945_));
 sky130_fd_sc_hd__clkbuf_1 _7995_ (.A(_3945_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _7996_ (.A0(\mem[20][21] ),
    .A1(_3791_),
    .S(_3944_),
    .X(_3946_));
 sky130_fd_sc_hd__clkbuf_1 _7997_ (.A(_3946_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _7998_ (.A0(\mem[20][22] ),
    .A1(_3793_),
    .S(_3944_),
    .X(_3947_));
 sky130_fd_sc_hd__clkbuf_1 _7999_ (.A(_3947_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _8000_ (.A0(\mem[20][23] ),
    .A1(_3795_),
    .S(_3944_),
    .X(_3948_));
 sky130_fd_sc_hd__clkbuf_1 _8001_ (.A(_3948_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _8002_ (.A0(\mem[20][24] ),
    .A1(_3797_),
    .S(_3944_),
    .X(_3949_));
 sky130_fd_sc_hd__clkbuf_1 _8003_ (.A(_3949_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _8004_ (.A0(\mem[20][25] ),
    .A1(_3799_),
    .S(_3944_),
    .X(_3950_));
 sky130_fd_sc_hd__clkbuf_1 _8005_ (.A(_3950_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _8006_ (.A0(\mem[20][26] ),
    .A1(_3801_),
    .S(_3944_),
    .X(_3951_));
 sky130_fd_sc_hd__clkbuf_1 _8007_ (.A(_3951_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _8008_ (.A0(\mem[20][27] ),
    .A1(_3803_),
    .S(_3944_),
    .X(_3952_));
 sky130_fd_sc_hd__clkbuf_1 _8009_ (.A(_3952_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _8010_ (.A0(\mem[20][28] ),
    .A1(_3805_),
    .S(_3944_),
    .X(_3953_));
 sky130_fd_sc_hd__clkbuf_1 _8011_ (.A(_3953_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _8012_ (.A0(\mem[20][29] ),
    .A1(_3807_),
    .S(_3944_),
    .X(_3954_));
 sky130_fd_sc_hd__clkbuf_1 _8013_ (.A(_3954_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _8014_ (.A0(\mem[20][30] ),
    .A1(_3809_),
    .S(_3921_),
    .X(_3955_));
 sky130_fd_sc_hd__clkbuf_1 _8015_ (.A(_3955_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _8016_ (.A0(\mem[20][31] ),
    .A1(_3811_),
    .S(_3921_),
    .X(_3956_));
 sky130_fd_sc_hd__clkbuf_1 _8017_ (.A(_3956_),
    .X(_0671_));
 sky130_fd_sc_hd__and3_4 _8018_ (.A(_3745_),
    .B(_3159_),
    .C(_3303_),
    .X(_3957_));
 sky130_fd_sc_hd__buf_6 _8019_ (.A(_3957_),
    .X(_3958_));
 sky130_fd_sc_hd__mux2_1 _8020_ (.A0(\mem[21][0] ),
    .A1(_3743_),
    .S(_3958_),
    .X(_3959_));
 sky130_fd_sc_hd__clkbuf_1 _8021_ (.A(_3959_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _8022_ (.A0(\mem[21][1] ),
    .A1(_3749_),
    .S(_3958_),
    .X(_3960_));
 sky130_fd_sc_hd__clkbuf_1 _8023_ (.A(_3960_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _8024_ (.A0(\mem[21][2] ),
    .A1(_3751_),
    .S(_3958_),
    .X(_3961_));
 sky130_fd_sc_hd__clkbuf_1 _8025_ (.A(_3961_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _8026_ (.A0(\mem[21][3] ),
    .A1(_3753_),
    .S(_3958_),
    .X(_3962_));
 sky130_fd_sc_hd__clkbuf_1 _8027_ (.A(_3962_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _8028_ (.A0(\mem[21][4] ),
    .A1(_3755_),
    .S(_3958_),
    .X(_3963_));
 sky130_fd_sc_hd__clkbuf_1 _8029_ (.A(_3963_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _8030_ (.A0(\mem[21][5] ),
    .A1(_3757_),
    .S(_3958_),
    .X(_3964_));
 sky130_fd_sc_hd__clkbuf_1 _8031_ (.A(_3964_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _8032_ (.A0(\mem[21][6] ),
    .A1(_3759_),
    .S(_3958_),
    .X(_3965_));
 sky130_fd_sc_hd__clkbuf_1 _8033_ (.A(_3965_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _8034_ (.A0(\mem[21][7] ),
    .A1(_3761_),
    .S(_3958_),
    .X(_3966_));
 sky130_fd_sc_hd__clkbuf_1 _8035_ (.A(_3966_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _8036_ (.A0(\mem[21][8] ),
    .A1(_3763_),
    .S(_3958_),
    .X(_3967_));
 sky130_fd_sc_hd__clkbuf_1 _8037_ (.A(_3967_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _8038_ (.A0(\mem[21][9] ),
    .A1(_3765_),
    .S(_3958_),
    .X(_3968_));
 sky130_fd_sc_hd__clkbuf_1 _8039_ (.A(_3968_),
    .X(_0681_));
 sky130_fd_sc_hd__buf_8 _8040_ (.A(_3957_),
    .X(_3969_));
 sky130_fd_sc_hd__mux2_1 _8041_ (.A0(\mem[21][10] ),
    .A1(_3767_),
    .S(_3969_),
    .X(_3970_));
 sky130_fd_sc_hd__clkbuf_1 _8042_ (.A(_3970_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _8043_ (.A0(\mem[21][11] ),
    .A1(_3770_),
    .S(_3969_),
    .X(_3971_));
 sky130_fd_sc_hd__clkbuf_1 _8044_ (.A(_3971_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _8045_ (.A0(\mem[21][12] ),
    .A1(_3772_),
    .S(_3969_),
    .X(_3972_));
 sky130_fd_sc_hd__clkbuf_1 _8046_ (.A(_3972_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _8047_ (.A0(\mem[21][13] ),
    .A1(_3774_),
    .S(_3969_),
    .X(_3973_));
 sky130_fd_sc_hd__clkbuf_1 _8048_ (.A(_3973_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _8049_ (.A0(\mem[21][14] ),
    .A1(_3776_),
    .S(_3969_),
    .X(_3974_));
 sky130_fd_sc_hd__clkbuf_1 _8050_ (.A(_3974_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _8051_ (.A0(\mem[21][15] ),
    .A1(_3778_),
    .S(_3969_),
    .X(_3975_));
 sky130_fd_sc_hd__clkbuf_1 _8052_ (.A(_3975_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _8053_ (.A0(\mem[21][16] ),
    .A1(_3780_),
    .S(_3969_),
    .X(_3976_));
 sky130_fd_sc_hd__clkbuf_1 _8054_ (.A(_3976_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _8055_ (.A0(\mem[21][17] ),
    .A1(_3782_),
    .S(_3969_),
    .X(_3977_));
 sky130_fd_sc_hd__clkbuf_1 _8056_ (.A(_3977_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _8057_ (.A0(\mem[21][18] ),
    .A1(_3784_),
    .S(_3969_),
    .X(_3978_));
 sky130_fd_sc_hd__clkbuf_1 _8058_ (.A(_3978_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _8059_ (.A0(\mem[21][19] ),
    .A1(_3786_),
    .S(_3969_),
    .X(_3979_));
 sky130_fd_sc_hd__clkbuf_1 _8060_ (.A(_3979_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_8 _8061_ (.A(_3957_),
    .X(_3980_));
 sky130_fd_sc_hd__mux2_1 _8062_ (.A0(\mem[21][20] ),
    .A1(_3788_),
    .S(_3980_),
    .X(_3981_));
 sky130_fd_sc_hd__clkbuf_1 _8063_ (.A(_3981_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _8064_ (.A0(\mem[21][21] ),
    .A1(_3791_),
    .S(_3980_),
    .X(_3982_));
 sky130_fd_sc_hd__clkbuf_1 _8065_ (.A(_3982_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _8066_ (.A0(\mem[21][22] ),
    .A1(_3793_),
    .S(_3980_),
    .X(_3983_));
 sky130_fd_sc_hd__clkbuf_1 _8067_ (.A(_3983_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _8068_ (.A0(\mem[21][23] ),
    .A1(_3795_),
    .S(_3980_),
    .X(_3984_));
 sky130_fd_sc_hd__clkbuf_1 _8069_ (.A(_3984_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _8070_ (.A0(\mem[21][24] ),
    .A1(_3797_),
    .S(_3980_),
    .X(_3985_));
 sky130_fd_sc_hd__clkbuf_1 _8071_ (.A(_3985_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _8072_ (.A0(\mem[21][25] ),
    .A1(_3799_),
    .S(_3980_),
    .X(_3986_));
 sky130_fd_sc_hd__clkbuf_1 _8073_ (.A(_3986_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _8074_ (.A0(\mem[21][26] ),
    .A1(_3801_),
    .S(_3980_),
    .X(_3987_));
 sky130_fd_sc_hd__clkbuf_1 _8075_ (.A(_3987_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _8076_ (.A0(\mem[21][27] ),
    .A1(_3803_),
    .S(_3980_),
    .X(_3988_));
 sky130_fd_sc_hd__clkbuf_1 _8077_ (.A(_3988_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _8078_ (.A0(\mem[21][28] ),
    .A1(_3805_),
    .S(_3980_),
    .X(_3989_));
 sky130_fd_sc_hd__clkbuf_1 _8079_ (.A(_3989_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _8080_ (.A0(\mem[21][29] ),
    .A1(_3807_),
    .S(_3980_),
    .X(_3990_));
 sky130_fd_sc_hd__clkbuf_1 _8081_ (.A(_3990_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _8082_ (.A0(\mem[21][30] ),
    .A1(_3809_),
    .S(_3957_),
    .X(_3991_));
 sky130_fd_sc_hd__clkbuf_1 _8083_ (.A(_3991_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _8084_ (.A0(\mem[21][31] ),
    .A1(_3811_),
    .S(_3957_),
    .X(_3992_));
 sky130_fd_sc_hd__clkbuf_1 _8085_ (.A(_3992_),
    .X(_0703_));
 sky130_fd_sc_hd__and3_2 _8086_ (.A(_3745_),
    .B(_3228_),
    .C(_3303_),
    .X(_3993_));
 sky130_fd_sc_hd__buf_4 _8087_ (.A(_3993_),
    .X(_3994_));
 sky130_fd_sc_hd__mux2_1 _8088_ (.A0(\mem[22][0] ),
    .A1(_3743_),
    .S(_3994_),
    .X(_3995_));
 sky130_fd_sc_hd__clkbuf_1 _8089_ (.A(_3995_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _8090_ (.A0(\mem[22][1] ),
    .A1(_3749_),
    .S(_3994_),
    .X(_3996_));
 sky130_fd_sc_hd__clkbuf_1 _8091_ (.A(_3996_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _8092_ (.A0(\mem[22][2] ),
    .A1(_3751_),
    .S(_3994_),
    .X(_3997_));
 sky130_fd_sc_hd__clkbuf_1 _8093_ (.A(_3997_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _8094_ (.A0(\mem[22][3] ),
    .A1(_3753_),
    .S(_3994_),
    .X(_3998_));
 sky130_fd_sc_hd__clkbuf_1 _8095_ (.A(_3998_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _8096_ (.A0(\mem[22][4] ),
    .A1(_3755_),
    .S(_3994_),
    .X(_3999_));
 sky130_fd_sc_hd__clkbuf_1 _8097_ (.A(_3999_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _8098_ (.A0(\mem[22][5] ),
    .A1(_3757_),
    .S(_3994_),
    .X(_4000_));
 sky130_fd_sc_hd__clkbuf_1 _8099_ (.A(_4000_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _8100_ (.A0(\mem[22][6] ),
    .A1(_3759_),
    .S(_3994_),
    .X(_4001_));
 sky130_fd_sc_hd__clkbuf_1 _8101_ (.A(_4001_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _8102_ (.A0(\mem[22][7] ),
    .A1(_3761_),
    .S(_3994_),
    .X(_4002_));
 sky130_fd_sc_hd__clkbuf_1 _8103_ (.A(_4002_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _8104_ (.A0(\mem[22][8] ),
    .A1(_3763_),
    .S(_3994_),
    .X(_4003_));
 sky130_fd_sc_hd__clkbuf_1 _8105_ (.A(_4003_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _8106_ (.A0(\mem[22][9] ),
    .A1(_3765_),
    .S(_3994_),
    .X(_4004_));
 sky130_fd_sc_hd__clkbuf_1 _8107_ (.A(_4004_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_6 _8108_ (.A(_3993_),
    .X(_4005_));
 sky130_fd_sc_hd__mux2_1 _8109_ (.A0(\mem[22][10] ),
    .A1(_3767_),
    .S(_4005_),
    .X(_4006_));
 sky130_fd_sc_hd__clkbuf_1 _8110_ (.A(_4006_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _8111_ (.A0(\mem[22][11] ),
    .A1(_3770_),
    .S(_4005_),
    .X(_4007_));
 sky130_fd_sc_hd__clkbuf_1 _8112_ (.A(_4007_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _8113_ (.A0(\mem[22][12] ),
    .A1(_3772_),
    .S(_4005_),
    .X(_4008_));
 sky130_fd_sc_hd__clkbuf_1 _8114_ (.A(_4008_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _8115_ (.A0(\mem[22][13] ),
    .A1(_3774_),
    .S(_4005_),
    .X(_4009_));
 sky130_fd_sc_hd__clkbuf_1 _8116_ (.A(_4009_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _8117_ (.A0(\mem[22][14] ),
    .A1(_3776_),
    .S(_4005_),
    .X(_4010_));
 sky130_fd_sc_hd__clkbuf_1 _8118_ (.A(_4010_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _8119_ (.A0(\mem[22][15] ),
    .A1(_3778_),
    .S(_4005_),
    .X(_4011_));
 sky130_fd_sc_hd__clkbuf_1 _8120_ (.A(_4011_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _8121_ (.A0(\mem[22][16] ),
    .A1(_3780_),
    .S(_4005_),
    .X(_4012_));
 sky130_fd_sc_hd__clkbuf_1 _8122_ (.A(_4012_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _8123_ (.A0(\mem[22][17] ),
    .A1(_3782_),
    .S(_4005_),
    .X(_4013_));
 sky130_fd_sc_hd__clkbuf_1 _8124_ (.A(_4013_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _8125_ (.A0(\mem[22][18] ),
    .A1(_3784_),
    .S(_4005_),
    .X(_4014_));
 sky130_fd_sc_hd__clkbuf_1 _8126_ (.A(_4014_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _8127_ (.A0(\mem[22][19] ),
    .A1(_3786_),
    .S(_4005_),
    .X(_4015_));
 sky130_fd_sc_hd__clkbuf_1 _8128_ (.A(_4015_),
    .X(_0723_));
 sky130_fd_sc_hd__buf_4 _8129_ (.A(_3993_),
    .X(_4016_));
 sky130_fd_sc_hd__mux2_1 _8130_ (.A0(\mem[22][20] ),
    .A1(_3788_),
    .S(_4016_),
    .X(_4017_));
 sky130_fd_sc_hd__clkbuf_1 _8131_ (.A(_4017_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _8132_ (.A0(\mem[22][21] ),
    .A1(_3791_),
    .S(_4016_),
    .X(_4018_));
 sky130_fd_sc_hd__clkbuf_1 _8133_ (.A(_4018_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _8134_ (.A0(\mem[22][22] ),
    .A1(_3793_),
    .S(_4016_),
    .X(_4019_));
 sky130_fd_sc_hd__clkbuf_1 _8135_ (.A(_4019_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _8136_ (.A0(\mem[22][23] ),
    .A1(_3795_),
    .S(_4016_),
    .X(_4020_));
 sky130_fd_sc_hd__clkbuf_1 _8137_ (.A(_4020_),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _8138_ (.A0(\mem[22][24] ),
    .A1(_3797_),
    .S(_4016_),
    .X(_4021_));
 sky130_fd_sc_hd__clkbuf_1 _8139_ (.A(_4021_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _8140_ (.A0(\mem[22][25] ),
    .A1(_3799_),
    .S(_4016_),
    .X(_4022_));
 sky130_fd_sc_hd__clkbuf_1 _8141_ (.A(_4022_),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _8142_ (.A0(\mem[22][26] ),
    .A1(_3801_),
    .S(_4016_),
    .X(_4023_));
 sky130_fd_sc_hd__clkbuf_1 _8143_ (.A(_4023_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _8144_ (.A0(\mem[22][27] ),
    .A1(_3803_),
    .S(_4016_),
    .X(_4024_));
 sky130_fd_sc_hd__clkbuf_1 _8145_ (.A(_4024_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _8146_ (.A0(\mem[22][28] ),
    .A1(_3805_),
    .S(_4016_),
    .X(_4025_));
 sky130_fd_sc_hd__clkbuf_1 _8147_ (.A(_4025_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _8148_ (.A0(\mem[22][29] ),
    .A1(_3807_),
    .S(_4016_),
    .X(_4026_));
 sky130_fd_sc_hd__clkbuf_1 _8149_ (.A(_4026_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _8150_ (.A0(\mem[22][30] ),
    .A1(_3809_),
    .S(_3993_),
    .X(_4027_));
 sky130_fd_sc_hd__clkbuf_1 _8151_ (.A(_4027_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _8152_ (.A0(\mem[22][31] ),
    .A1(_3811_),
    .S(_3993_),
    .X(_4028_));
 sky130_fd_sc_hd__clkbuf_1 _8153_ (.A(_4028_),
    .X(_0735_));
 sky130_fd_sc_hd__or3_4 _8154_ (.A(_3087_),
    .B(_3088_),
    .C(_3341_),
    .X(_4029_));
 sky130_fd_sc_hd__buf_4 _8155_ (.A(_4029_),
    .X(_4030_));
 sky130_fd_sc_hd__mux2_1 _8156_ (.A0(_3086_),
    .A1(\mem[23][0] ),
    .S(_4030_),
    .X(_4031_));
 sky130_fd_sc_hd__clkbuf_1 _8157_ (.A(_4031_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _8158_ (.A0(_3093_),
    .A1(\mem[23][1] ),
    .S(_4030_),
    .X(_4032_));
 sky130_fd_sc_hd__clkbuf_1 _8159_ (.A(_4032_),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _8160_ (.A0(_3095_),
    .A1(\mem[23][2] ),
    .S(_4030_),
    .X(_4033_));
 sky130_fd_sc_hd__clkbuf_1 _8161_ (.A(_4033_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _8162_ (.A0(_3097_),
    .A1(\mem[23][3] ),
    .S(_4030_),
    .X(_4034_));
 sky130_fd_sc_hd__clkbuf_1 _8163_ (.A(_4034_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _8164_ (.A0(_3099_),
    .A1(\mem[23][4] ),
    .S(_4030_),
    .X(_4035_));
 sky130_fd_sc_hd__clkbuf_1 _8165_ (.A(_4035_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _8166_ (.A0(_3101_),
    .A1(\mem[23][5] ),
    .S(_4030_),
    .X(_4036_));
 sky130_fd_sc_hd__clkbuf_1 _8167_ (.A(_4036_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _8168_ (.A0(_3103_),
    .A1(\mem[23][6] ),
    .S(_4030_),
    .X(_4037_));
 sky130_fd_sc_hd__clkbuf_1 _8169_ (.A(_4037_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _8170_ (.A0(_3105_),
    .A1(\mem[23][7] ),
    .S(_4030_),
    .X(_4038_));
 sky130_fd_sc_hd__clkbuf_1 _8171_ (.A(_4038_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _8172_ (.A0(_3107_),
    .A1(\mem[23][8] ),
    .S(_4030_),
    .X(_4039_));
 sky130_fd_sc_hd__clkbuf_1 _8173_ (.A(_4039_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _8174_ (.A0(_3109_),
    .A1(\mem[23][9] ),
    .S(_4030_),
    .X(_4040_));
 sky130_fd_sc_hd__clkbuf_1 _8175_ (.A(_4040_),
    .X(_0745_));
 sky130_fd_sc_hd__buf_6 _8176_ (.A(_4029_),
    .X(_4041_));
 sky130_fd_sc_hd__mux2_1 _8177_ (.A0(_3111_),
    .A1(\mem[23][10] ),
    .S(_4041_),
    .X(_4042_));
 sky130_fd_sc_hd__clkbuf_1 _8178_ (.A(_4042_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _8179_ (.A0(_3114_),
    .A1(\mem[23][11] ),
    .S(_4041_),
    .X(_4043_));
 sky130_fd_sc_hd__clkbuf_1 _8180_ (.A(_4043_),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _8181_ (.A0(_3116_),
    .A1(\mem[23][12] ),
    .S(_4041_),
    .X(_4044_));
 sky130_fd_sc_hd__clkbuf_1 _8182_ (.A(_4044_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _8183_ (.A0(_3118_),
    .A1(\mem[23][13] ),
    .S(_4041_),
    .X(_4045_));
 sky130_fd_sc_hd__clkbuf_1 _8184_ (.A(_4045_),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _8185_ (.A0(_3120_),
    .A1(\mem[23][14] ),
    .S(_4041_),
    .X(_4046_));
 sky130_fd_sc_hd__clkbuf_1 _8186_ (.A(_4046_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _8187_ (.A0(_3122_),
    .A1(\mem[23][15] ),
    .S(_4041_),
    .X(_4047_));
 sky130_fd_sc_hd__clkbuf_1 _8188_ (.A(_4047_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _8189_ (.A0(_3124_),
    .A1(\mem[23][16] ),
    .S(_4041_),
    .X(_4048_));
 sky130_fd_sc_hd__clkbuf_1 _8190_ (.A(_4048_),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _8191_ (.A0(_3126_),
    .A1(\mem[23][17] ),
    .S(_4041_),
    .X(_4049_));
 sky130_fd_sc_hd__clkbuf_1 _8192_ (.A(_4049_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _8193_ (.A0(_3128_),
    .A1(\mem[23][18] ),
    .S(_4041_),
    .X(_4050_));
 sky130_fd_sc_hd__clkbuf_1 _8194_ (.A(_4050_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _8195_ (.A0(_3130_),
    .A1(\mem[23][19] ),
    .S(_4041_),
    .X(_4051_));
 sky130_fd_sc_hd__clkbuf_1 _8196_ (.A(_4051_),
    .X(_0755_));
 sky130_fd_sc_hd__buf_4 _8197_ (.A(_4029_),
    .X(_4052_));
 sky130_fd_sc_hd__mux2_1 _8198_ (.A0(_3132_),
    .A1(\mem[23][20] ),
    .S(_4052_),
    .X(_4053_));
 sky130_fd_sc_hd__clkbuf_1 _8199_ (.A(_4053_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _8200_ (.A0(_3135_),
    .A1(\mem[23][21] ),
    .S(_4052_),
    .X(_4054_));
 sky130_fd_sc_hd__clkbuf_1 _8201_ (.A(_4054_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _8202_ (.A0(_3137_),
    .A1(\mem[23][22] ),
    .S(_4052_),
    .X(_4055_));
 sky130_fd_sc_hd__clkbuf_1 _8203_ (.A(_4055_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _8204_ (.A0(_3139_),
    .A1(\mem[23][23] ),
    .S(_4052_),
    .X(_4056_));
 sky130_fd_sc_hd__clkbuf_1 _8205_ (.A(_4056_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _8206_ (.A0(_3141_),
    .A1(\mem[23][24] ),
    .S(_4052_),
    .X(_4057_));
 sky130_fd_sc_hd__clkbuf_1 _8207_ (.A(_4057_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _8208_ (.A0(_3143_),
    .A1(\mem[23][25] ),
    .S(_4052_),
    .X(_4058_));
 sky130_fd_sc_hd__clkbuf_1 _8209_ (.A(_4058_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _8210_ (.A0(_3145_),
    .A1(\mem[23][26] ),
    .S(_4052_),
    .X(_4059_));
 sky130_fd_sc_hd__clkbuf_1 _8211_ (.A(_4059_),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_1 _8212_ (.A0(_3147_),
    .A1(\mem[23][27] ),
    .S(_4052_),
    .X(_4060_));
 sky130_fd_sc_hd__clkbuf_1 _8213_ (.A(_4060_),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _8214_ (.A0(_3149_),
    .A1(\mem[23][28] ),
    .S(_4052_),
    .X(_4061_));
 sky130_fd_sc_hd__clkbuf_1 _8215_ (.A(_4061_),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _8216_ (.A0(_3151_),
    .A1(\mem[23][29] ),
    .S(_4052_),
    .X(_4062_));
 sky130_fd_sc_hd__clkbuf_1 _8217_ (.A(_4062_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _8218_ (.A0(_3153_),
    .A1(\mem[23][30] ),
    .S(_4029_),
    .X(_4063_));
 sky130_fd_sc_hd__clkbuf_1 _8219_ (.A(_4063_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _8220_ (.A0(_3155_),
    .A1(\mem[23][31] ),
    .S(_4029_),
    .X(_4064_));
 sky130_fd_sc_hd__clkbuf_1 _8221_ (.A(_4064_),
    .X(_0767_));
 sky130_fd_sc_hd__and3_2 _8222_ (.A(_3745_),
    .B(_3302_),
    .C(_3452_),
    .X(_4065_));
 sky130_fd_sc_hd__buf_6 _8223_ (.A(_4065_),
    .X(_4066_));
 sky130_fd_sc_hd__mux2_1 _8224_ (.A0(\mem[24][0] ),
    .A1(_3743_),
    .S(_4066_),
    .X(_4067_));
 sky130_fd_sc_hd__clkbuf_1 _8225_ (.A(_4067_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _8226_ (.A0(\mem[24][1] ),
    .A1(_3749_),
    .S(_4066_),
    .X(_4068_));
 sky130_fd_sc_hd__clkbuf_1 _8227_ (.A(_4068_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _8228_ (.A0(\mem[24][2] ),
    .A1(_3751_),
    .S(_4066_),
    .X(_4069_));
 sky130_fd_sc_hd__clkbuf_1 _8229_ (.A(_4069_),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _8230_ (.A0(\mem[24][3] ),
    .A1(_3753_),
    .S(_4066_),
    .X(_4070_));
 sky130_fd_sc_hd__clkbuf_1 _8231_ (.A(_4070_),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _8232_ (.A0(\mem[24][4] ),
    .A1(_3755_),
    .S(_4066_),
    .X(_4071_));
 sky130_fd_sc_hd__clkbuf_1 _8233_ (.A(_4071_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _8234_ (.A0(\mem[24][5] ),
    .A1(_3757_),
    .S(_4066_),
    .X(_4072_));
 sky130_fd_sc_hd__clkbuf_1 _8235_ (.A(_4072_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _8236_ (.A0(\mem[24][6] ),
    .A1(_3759_),
    .S(_4066_),
    .X(_4073_));
 sky130_fd_sc_hd__clkbuf_1 _8237_ (.A(_4073_),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _8238_ (.A0(\mem[24][7] ),
    .A1(_3761_),
    .S(_4066_),
    .X(_4074_));
 sky130_fd_sc_hd__clkbuf_1 _8239_ (.A(_4074_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _8240_ (.A0(\mem[24][8] ),
    .A1(_3763_),
    .S(_4066_),
    .X(_4075_));
 sky130_fd_sc_hd__clkbuf_1 _8241_ (.A(_4075_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _8242_ (.A0(\mem[24][9] ),
    .A1(_3765_),
    .S(_4066_),
    .X(_4076_));
 sky130_fd_sc_hd__clkbuf_1 _8243_ (.A(_4076_),
    .X(_0777_));
 sky130_fd_sc_hd__clkbuf_8 _8244_ (.A(_4065_),
    .X(_4077_));
 sky130_fd_sc_hd__mux2_1 _8245_ (.A0(\mem[24][10] ),
    .A1(_3767_),
    .S(_4077_),
    .X(_4078_));
 sky130_fd_sc_hd__clkbuf_1 _8246_ (.A(_4078_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _8247_ (.A0(\mem[24][11] ),
    .A1(_3770_),
    .S(_4077_),
    .X(_4079_));
 sky130_fd_sc_hd__clkbuf_1 _8248_ (.A(_4079_),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _8249_ (.A0(\mem[24][12] ),
    .A1(_3772_),
    .S(_4077_),
    .X(_4080_));
 sky130_fd_sc_hd__clkbuf_1 _8250_ (.A(_4080_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _8251_ (.A0(\mem[24][13] ),
    .A1(_3774_),
    .S(_4077_),
    .X(_4081_));
 sky130_fd_sc_hd__clkbuf_1 _8252_ (.A(_4081_),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _8253_ (.A0(\mem[24][14] ),
    .A1(_3776_),
    .S(_4077_),
    .X(_4082_));
 sky130_fd_sc_hd__clkbuf_1 _8254_ (.A(_4082_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _8255_ (.A0(\mem[24][15] ),
    .A1(_3778_),
    .S(_4077_),
    .X(_4083_));
 sky130_fd_sc_hd__clkbuf_1 _8256_ (.A(_4083_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _8257_ (.A0(\mem[24][16] ),
    .A1(_3780_),
    .S(_4077_),
    .X(_4084_));
 sky130_fd_sc_hd__clkbuf_1 _8258_ (.A(_4084_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _8259_ (.A0(\mem[24][17] ),
    .A1(_3782_),
    .S(_4077_),
    .X(_4085_));
 sky130_fd_sc_hd__clkbuf_1 _8260_ (.A(_4085_),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _8261_ (.A0(\mem[24][18] ),
    .A1(_3784_),
    .S(_4077_),
    .X(_4086_));
 sky130_fd_sc_hd__clkbuf_1 _8262_ (.A(_4086_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _8263_ (.A0(\mem[24][19] ),
    .A1(_3786_),
    .S(_4077_),
    .X(_4087_));
 sky130_fd_sc_hd__clkbuf_1 _8264_ (.A(_4087_),
    .X(_0787_));
 sky130_fd_sc_hd__buf_4 _8265_ (.A(_4065_),
    .X(_4088_));
 sky130_fd_sc_hd__mux2_1 _8266_ (.A0(\mem[24][20] ),
    .A1(_3788_),
    .S(_4088_),
    .X(_4089_));
 sky130_fd_sc_hd__clkbuf_1 _8267_ (.A(_4089_),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _8268_ (.A0(\mem[24][21] ),
    .A1(_3791_),
    .S(_4088_),
    .X(_4090_));
 sky130_fd_sc_hd__clkbuf_1 _8269_ (.A(_4090_),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _8270_ (.A0(\mem[24][22] ),
    .A1(_3793_),
    .S(_4088_),
    .X(_4091_));
 sky130_fd_sc_hd__clkbuf_1 _8271_ (.A(_4091_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _8272_ (.A0(\mem[24][23] ),
    .A1(_3795_),
    .S(_4088_),
    .X(_4092_));
 sky130_fd_sc_hd__clkbuf_1 _8273_ (.A(_4092_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _8274_ (.A0(\mem[24][24] ),
    .A1(_3797_),
    .S(_4088_),
    .X(_4093_));
 sky130_fd_sc_hd__clkbuf_1 _8275_ (.A(_4093_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _8276_ (.A0(\mem[24][25] ),
    .A1(_3799_),
    .S(_4088_),
    .X(_4094_));
 sky130_fd_sc_hd__clkbuf_1 _8277_ (.A(_4094_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _8278_ (.A0(\mem[24][26] ),
    .A1(_3801_),
    .S(_4088_),
    .X(_4095_));
 sky130_fd_sc_hd__clkbuf_1 _8279_ (.A(_4095_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _8280_ (.A0(\mem[24][27] ),
    .A1(_3803_),
    .S(_4088_),
    .X(_4096_));
 sky130_fd_sc_hd__clkbuf_1 _8281_ (.A(_4096_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _8282_ (.A0(\mem[24][28] ),
    .A1(_3805_),
    .S(_4088_),
    .X(_4097_));
 sky130_fd_sc_hd__clkbuf_1 _8283_ (.A(_4097_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _8284_ (.A0(\mem[24][29] ),
    .A1(_3807_),
    .S(_4088_),
    .X(_4098_));
 sky130_fd_sc_hd__clkbuf_1 _8285_ (.A(_4098_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _8286_ (.A0(\mem[24][30] ),
    .A1(_3809_),
    .S(_4065_),
    .X(_4099_));
 sky130_fd_sc_hd__clkbuf_1 _8287_ (.A(_4099_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _8288_ (.A0(\mem[24][31] ),
    .A1(_3811_),
    .S(_4065_),
    .X(_4100_));
 sky130_fd_sc_hd__clkbuf_1 _8289_ (.A(_4100_),
    .X(_0799_));
 sky130_fd_sc_hd__and3_4 _8290_ (.A(_3745_),
    .B(_3159_),
    .C(_3452_),
    .X(_4101_));
 sky130_fd_sc_hd__buf_6 _8291_ (.A(_4101_),
    .X(_4102_));
 sky130_fd_sc_hd__mux2_1 _8292_ (.A0(\mem[25][0] ),
    .A1(_3743_),
    .S(_4102_),
    .X(_4103_));
 sky130_fd_sc_hd__clkbuf_1 _8293_ (.A(_4103_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _8294_ (.A0(\mem[25][1] ),
    .A1(_3749_),
    .S(_4102_),
    .X(_4104_));
 sky130_fd_sc_hd__clkbuf_1 _8295_ (.A(_4104_),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _8296_ (.A0(\mem[25][2] ),
    .A1(_3751_),
    .S(_4102_),
    .X(_4105_));
 sky130_fd_sc_hd__clkbuf_1 _8297_ (.A(_4105_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _8298_ (.A0(\mem[25][3] ),
    .A1(_3753_),
    .S(_4102_),
    .X(_4106_));
 sky130_fd_sc_hd__clkbuf_1 _8299_ (.A(_4106_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _8300_ (.A0(\mem[25][4] ),
    .A1(_3755_),
    .S(_4102_),
    .X(_4107_));
 sky130_fd_sc_hd__clkbuf_1 _8301_ (.A(_4107_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _8302_ (.A0(\mem[25][5] ),
    .A1(_3757_),
    .S(_4102_),
    .X(_4108_));
 sky130_fd_sc_hd__clkbuf_1 _8303_ (.A(_4108_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _8304_ (.A0(\mem[25][6] ),
    .A1(_3759_),
    .S(_4102_),
    .X(_4109_));
 sky130_fd_sc_hd__clkbuf_1 _8305_ (.A(_4109_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _8306_ (.A0(\mem[25][7] ),
    .A1(_3761_),
    .S(_4102_),
    .X(_4110_));
 sky130_fd_sc_hd__clkbuf_1 _8307_ (.A(_4110_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _8308_ (.A0(\mem[25][8] ),
    .A1(_3763_),
    .S(_4102_),
    .X(_4111_));
 sky130_fd_sc_hd__clkbuf_1 _8309_ (.A(_4111_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _8310_ (.A0(\mem[25][9] ),
    .A1(_3765_),
    .S(_4102_),
    .X(_4112_));
 sky130_fd_sc_hd__clkbuf_1 _8311_ (.A(_4112_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_6 _8312_ (.A(_4101_),
    .X(_4113_));
 sky130_fd_sc_hd__mux2_1 _8313_ (.A0(\mem[25][10] ),
    .A1(_3767_),
    .S(_4113_),
    .X(_4114_));
 sky130_fd_sc_hd__clkbuf_1 _8314_ (.A(_4114_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _8315_ (.A0(\mem[25][11] ),
    .A1(_3770_),
    .S(_4113_),
    .X(_4115_));
 sky130_fd_sc_hd__clkbuf_1 _8316_ (.A(_4115_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _8317_ (.A0(\mem[25][12] ),
    .A1(_3772_),
    .S(_4113_),
    .X(_4116_));
 sky130_fd_sc_hd__clkbuf_1 _8318_ (.A(_4116_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _8319_ (.A0(\mem[25][13] ),
    .A1(_3774_),
    .S(_4113_),
    .X(_4117_));
 sky130_fd_sc_hd__clkbuf_1 _8320_ (.A(_4117_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _8321_ (.A0(\mem[25][14] ),
    .A1(_3776_),
    .S(_4113_),
    .X(_4118_));
 sky130_fd_sc_hd__clkbuf_1 _8322_ (.A(_4118_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _8323_ (.A0(\mem[25][15] ),
    .A1(_3778_),
    .S(_4113_),
    .X(_4119_));
 sky130_fd_sc_hd__clkbuf_1 _8324_ (.A(_4119_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _8325_ (.A0(\mem[25][16] ),
    .A1(_3780_),
    .S(_4113_),
    .X(_4120_));
 sky130_fd_sc_hd__clkbuf_1 _8326_ (.A(_4120_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _8327_ (.A0(\mem[25][17] ),
    .A1(_3782_),
    .S(_4113_),
    .X(_4121_));
 sky130_fd_sc_hd__clkbuf_1 _8328_ (.A(_4121_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _8329_ (.A0(\mem[25][18] ),
    .A1(_3784_),
    .S(_4113_),
    .X(_4122_));
 sky130_fd_sc_hd__clkbuf_1 _8330_ (.A(_4122_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _8331_ (.A0(\mem[25][19] ),
    .A1(_3786_),
    .S(_4113_),
    .X(_4123_));
 sky130_fd_sc_hd__clkbuf_1 _8332_ (.A(_4123_),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _8333_ (.A(_4101_),
    .X(_4124_));
 sky130_fd_sc_hd__mux2_1 _8334_ (.A0(\mem[25][20] ),
    .A1(_3788_),
    .S(_4124_),
    .X(_4125_));
 sky130_fd_sc_hd__clkbuf_1 _8335_ (.A(_4125_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _8336_ (.A0(\mem[25][21] ),
    .A1(_3791_),
    .S(_4124_),
    .X(_4126_));
 sky130_fd_sc_hd__clkbuf_1 _8337_ (.A(_4126_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _8338_ (.A0(\mem[25][22] ),
    .A1(_3793_),
    .S(_4124_),
    .X(_4127_));
 sky130_fd_sc_hd__clkbuf_1 _8339_ (.A(_4127_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _8340_ (.A0(\mem[25][23] ),
    .A1(_3795_),
    .S(_4124_),
    .X(_4128_));
 sky130_fd_sc_hd__clkbuf_1 _8341_ (.A(_4128_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _8342_ (.A0(\mem[25][24] ),
    .A1(_3797_),
    .S(_4124_),
    .X(_4129_));
 sky130_fd_sc_hd__clkbuf_1 _8343_ (.A(_4129_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _8344_ (.A0(\mem[25][25] ),
    .A1(_3799_),
    .S(_4124_),
    .X(_4130_));
 sky130_fd_sc_hd__clkbuf_1 _8345_ (.A(_4130_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _8346_ (.A0(\mem[25][26] ),
    .A1(_3801_),
    .S(_4124_),
    .X(_4131_));
 sky130_fd_sc_hd__clkbuf_1 _8347_ (.A(_4131_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _8348_ (.A0(\mem[25][27] ),
    .A1(_3803_),
    .S(_4124_),
    .X(_4132_));
 sky130_fd_sc_hd__clkbuf_1 _8349_ (.A(_4132_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _8350_ (.A0(\mem[25][28] ),
    .A1(_3805_),
    .S(_4124_),
    .X(_4133_));
 sky130_fd_sc_hd__clkbuf_1 _8351_ (.A(_4133_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _8352_ (.A0(\mem[25][29] ),
    .A1(_3807_),
    .S(_4124_),
    .X(_4134_));
 sky130_fd_sc_hd__clkbuf_1 _8353_ (.A(_4134_),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _8354_ (.A0(\mem[25][30] ),
    .A1(_3809_),
    .S(_4101_),
    .X(_4135_));
 sky130_fd_sc_hd__clkbuf_1 _8355_ (.A(_4135_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _8356_ (.A0(\mem[25][31] ),
    .A1(_3811_),
    .S(_4101_),
    .X(_4136_));
 sky130_fd_sc_hd__clkbuf_1 _8357_ (.A(_4136_),
    .X(_0831_));
 sky130_fd_sc_hd__and3_4 _8358_ (.A(_3745_),
    .B(_3228_),
    .C(_3452_),
    .X(_4137_));
 sky130_fd_sc_hd__buf_6 _8359_ (.A(_4137_),
    .X(_4138_));
 sky130_fd_sc_hd__mux2_1 _8360_ (.A0(\mem[26][0] ),
    .A1(_3743_),
    .S(_4138_),
    .X(_4139_));
 sky130_fd_sc_hd__clkbuf_1 _8361_ (.A(_4139_),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _8362_ (.A0(\mem[26][1] ),
    .A1(_3749_),
    .S(_4138_),
    .X(_4140_));
 sky130_fd_sc_hd__clkbuf_1 _8363_ (.A(_4140_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _8364_ (.A0(\mem[26][2] ),
    .A1(_3751_),
    .S(_4138_),
    .X(_4141_));
 sky130_fd_sc_hd__clkbuf_1 _8365_ (.A(_4141_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _8366_ (.A0(\mem[26][3] ),
    .A1(_3753_),
    .S(_4138_),
    .X(_4142_));
 sky130_fd_sc_hd__clkbuf_1 _8367_ (.A(_4142_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _8368_ (.A0(\mem[26][4] ),
    .A1(_3755_),
    .S(_4138_),
    .X(_4143_));
 sky130_fd_sc_hd__clkbuf_1 _8369_ (.A(_4143_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _8370_ (.A0(\mem[26][5] ),
    .A1(_3757_),
    .S(_4138_),
    .X(_4144_));
 sky130_fd_sc_hd__clkbuf_1 _8371_ (.A(_4144_),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _8372_ (.A0(\mem[26][6] ),
    .A1(_3759_),
    .S(_4138_),
    .X(_4145_));
 sky130_fd_sc_hd__clkbuf_1 _8373_ (.A(_4145_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _8374_ (.A0(\mem[26][7] ),
    .A1(_3761_),
    .S(_4138_),
    .X(_4146_));
 sky130_fd_sc_hd__clkbuf_1 _8375_ (.A(_4146_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _8376_ (.A0(\mem[26][8] ),
    .A1(_3763_),
    .S(_4138_),
    .X(_4147_));
 sky130_fd_sc_hd__clkbuf_1 _8377_ (.A(_4147_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _8378_ (.A0(\mem[26][9] ),
    .A1(_3765_),
    .S(_4138_),
    .X(_4148_));
 sky130_fd_sc_hd__clkbuf_1 _8379_ (.A(_4148_),
    .X(_0841_));
 sky130_fd_sc_hd__buf_6 _8380_ (.A(_4137_),
    .X(_4149_));
 sky130_fd_sc_hd__mux2_1 _8381_ (.A0(\mem[26][10] ),
    .A1(_3767_),
    .S(_4149_),
    .X(_4150_));
 sky130_fd_sc_hd__clkbuf_1 _8382_ (.A(_4150_),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _8383_ (.A0(\mem[26][11] ),
    .A1(_3770_),
    .S(_4149_),
    .X(_4151_));
 sky130_fd_sc_hd__clkbuf_1 _8384_ (.A(_4151_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _8385_ (.A0(\mem[26][12] ),
    .A1(_3772_),
    .S(_4149_),
    .X(_4152_));
 sky130_fd_sc_hd__clkbuf_1 _8386_ (.A(_4152_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _8387_ (.A0(\mem[26][13] ),
    .A1(_3774_),
    .S(_4149_),
    .X(_4153_));
 sky130_fd_sc_hd__clkbuf_1 _8388_ (.A(_4153_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _8389_ (.A0(\mem[26][14] ),
    .A1(_3776_),
    .S(_4149_),
    .X(_4154_));
 sky130_fd_sc_hd__clkbuf_1 _8390_ (.A(_4154_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _8391_ (.A0(\mem[26][15] ),
    .A1(_3778_),
    .S(_4149_),
    .X(_4155_));
 sky130_fd_sc_hd__clkbuf_1 _8392_ (.A(_4155_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _8393_ (.A0(\mem[26][16] ),
    .A1(_3780_),
    .S(_4149_),
    .X(_4156_));
 sky130_fd_sc_hd__clkbuf_1 _8394_ (.A(_4156_),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _8395_ (.A0(\mem[26][17] ),
    .A1(_3782_),
    .S(_4149_),
    .X(_4157_));
 sky130_fd_sc_hd__clkbuf_1 _8396_ (.A(_4157_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _8397_ (.A0(\mem[26][18] ),
    .A1(_3784_),
    .S(_4149_),
    .X(_4158_));
 sky130_fd_sc_hd__clkbuf_1 _8398_ (.A(_4158_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _8399_ (.A0(\mem[26][19] ),
    .A1(_3786_),
    .S(_4149_),
    .X(_4159_));
 sky130_fd_sc_hd__clkbuf_1 _8400_ (.A(_4159_),
    .X(_0851_));
 sky130_fd_sc_hd__buf_4 _8401_ (.A(_4137_),
    .X(_4160_));
 sky130_fd_sc_hd__mux2_1 _8402_ (.A0(\mem[26][20] ),
    .A1(_3788_),
    .S(_4160_),
    .X(_4161_));
 sky130_fd_sc_hd__clkbuf_1 _8403_ (.A(_4161_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _8404_ (.A0(\mem[26][21] ),
    .A1(_3791_),
    .S(_4160_),
    .X(_4162_));
 sky130_fd_sc_hd__clkbuf_1 _8405_ (.A(_4162_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _8406_ (.A0(\mem[26][22] ),
    .A1(_3793_),
    .S(_4160_),
    .X(_4163_));
 sky130_fd_sc_hd__clkbuf_1 _8407_ (.A(_4163_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _8408_ (.A0(\mem[26][23] ),
    .A1(_3795_),
    .S(_4160_),
    .X(_4164_));
 sky130_fd_sc_hd__clkbuf_1 _8409_ (.A(_4164_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _8410_ (.A0(\mem[26][24] ),
    .A1(_3797_),
    .S(_4160_),
    .X(_4165_));
 sky130_fd_sc_hd__clkbuf_1 _8411_ (.A(_4165_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _8412_ (.A0(\mem[26][25] ),
    .A1(_3799_),
    .S(_4160_),
    .X(_4166_));
 sky130_fd_sc_hd__clkbuf_1 _8413_ (.A(_4166_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _8414_ (.A0(\mem[26][26] ),
    .A1(_3801_),
    .S(_4160_),
    .X(_4167_));
 sky130_fd_sc_hd__clkbuf_1 _8415_ (.A(_4167_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _8416_ (.A0(\mem[26][27] ),
    .A1(_3803_),
    .S(_4160_),
    .X(_4168_));
 sky130_fd_sc_hd__clkbuf_1 _8417_ (.A(_4168_),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _8418_ (.A0(\mem[26][28] ),
    .A1(_3805_),
    .S(_4160_),
    .X(_4169_));
 sky130_fd_sc_hd__clkbuf_1 _8419_ (.A(_4169_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _8420_ (.A0(\mem[26][29] ),
    .A1(_3807_),
    .S(_4160_),
    .X(_4170_));
 sky130_fd_sc_hd__clkbuf_1 _8421_ (.A(_4170_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _8422_ (.A0(\mem[26][30] ),
    .A1(_3809_),
    .S(_4137_),
    .X(_4171_));
 sky130_fd_sc_hd__clkbuf_1 _8423_ (.A(_4171_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _8424_ (.A0(\mem[26][31] ),
    .A1(_3811_),
    .S(_4137_),
    .X(_4172_));
 sky130_fd_sc_hd__clkbuf_1 _8425_ (.A(_4172_),
    .X(_0863_));
 sky130_fd_sc_hd__or3_4 _8426_ (.A(_3087_),
    .B(_3088_),
    .C(_3489_),
    .X(_4173_));
 sky130_fd_sc_hd__buf_6 _8427_ (.A(_4173_),
    .X(_4174_));
 sky130_fd_sc_hd__mux2_1 _8428_ (.A0(_3086_),
    .A1(\mem[27][0] ),
    .S(_4174_),
    .X(_4175_));
 sky130_fd_sc_hd__clkbuf_1 _8429_ (.A(_4175_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _8430_ (.A0(_3093_),
    .A1(\mem[27][1] ),
    .S(_4174_),
    .X(_4176_));
 sky130_fd_sc_hd__clkbuf_1 _8431_ (.A(_4176_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _8432_ (.A0(_3095_),
    .A1(\mem[27][2] ),
    .S(_4174_),
    .X(_4177_));
 sky130_fd_sc_hd__clkbuf_1 _8433_ (.A(_4177_),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _8434_ (.A0(_3097_),
    .A1(\mem[27][3] ),
    .S(_4174_),
    .X(_4178_));
 sky130_fd_sc_hd__clkbuf_1 _8435_ (.A(_4178_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _8436_ (.A0(_3099_),
    .A1(\mem[27][4] ),
    .S(_4174_),
    .X(_4179_));
 sky130_fd_sc_hd__clkbuf_1 _8437_ (.A(_4179_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _8438_ (.A0(_3101_),
    .A1(\mem[27][5] ),
    .S(_4174_),
    .X(_4180_));
 sky130_fd_sc_hd__clkbuf_1 _8439_ (.A(_4180_),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _8440_ (.A0(_3103_),
    .A1(\mem[27][6] ),
    .S(_4174_),
    .X(_4181_));
 sky130_fd_sc_hd__clkbuf_1 _8441_ (.A(_4181_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _8442_ (.A0(_3105_),
    .A1(\mem[27][7] ),
    .S(_4174_),
    .X(_4182_));
 sky130_fd_sc_hd__clkbuf_1 _8443_ (.A(_4182_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _8444_ (.A0(_3107_),
    .A1(\mem[27][8] ),
    .S(_4174_),
    .X(_4183_));
 sky130_fd_sc_hd__clkbuf_1 _8445_ (.A(_4183_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _8446_ (.A0(_3109_),
    .A1(\mem[27][9] ),
    .S(_4174_),
    .X(_4184_));
 sky130_fd_sc_hd__clkbuf_1 _8447_ (.A(_4184_),
    .X(_0873_));
 sky130_fd_sc_hd__buf_6 _8448_ (.A(_4173_),
    .X(_4185_));
 sky130_fd_sc_hd__mux2_1 _8449_ (.A0(_3111_),
    .A1(\mem[27][10] ),
    .S(_4185_),
    .X(_4186_));
 sky130_fd_sc_hd__clkbuf_1 _8450_ (.A(_4186_),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _8451_ (.A0(_3114_),
    .A1(\mem[27][11] ),
    .S(_4185_),
    .X(_4187_));
 sky130_fd_sc_hd__clkbuf_1 _8452_ (.A(_4187_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _8453_ (.A0(_3116_),
    .A1(\mem[27][12] ),
    .S(_4185_),
    .X(_4188_));
 sky130_fd_sc_hd__clkbuf_1 _8454_ (.A(_4188_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _8455_ (.A0(_3118_),
    .A1(\mem[27][13] ),
    .S(_4185_),
    .X(_4189_));
 sky130_fd_sc_hd__clkbuf_1 _8456_ (.A(_4189_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _8457_ (.A0(_3120_),
    .A1(\mem[27][14] ),
    .S(_4185_),
    .X(_4190_));
 sky130_fd_sc_hd__clkbuf_1 _8458_ (.A(_4190_),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _8459_ (.A0(_3122_),
    .A1(\mem[27][15] ),
    .S(_4185_),
    .X(_4191_));
 sky130_fd_sc_hd__clkbuf_1 _8460_ (.A(_4191_),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_1 _8461_ (.A0(_3124_),
    .A1(\mem[27][16] ),
    .S(_4185_),
    .X(_4192_));
 sky130_fd_sc_hd__clkbuf_1 _8462_ (.A(_4192_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _8463_ (.A0(_3126_),
    .A1(\mem[27][17] ),
    .S(_4185_),
    .X(_4193_));
 sky130_fd_sc_hd__clkbuf_1 _8464_ (.A(_4193_),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _8465_ (.A0(_3128_),
    .A1(\mem[27][18] ),
    .S(_4185_),
    .X(_4194_));
 sky130_fd_sc_hd__clkbuf_1 _8466_ (.A(_4194_),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _8467_ (.A0(_3130_),
    .A1(\mem[27][19] ),
    .S(_4185_),
    .X(_4195_));
 sky130_fd_sc_hd__clkbuf_1 _8468_ (.A(_4195_),
    .X(_0883_));
 sky130_fd_sc_hd__buf_4 _8469_ (.A(_4173_),
    .X(_4196_));
 sky130_fd_sc_hd__mux2_1 _8470_ (.A0(_3132_),
    .A1(\mem[27][20] ),
    .S(_4196_),
    .X(_4197_));
 sky130_fd_sc_hd__clkbuf_1 _8471_ (.A(_4197_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _8472_ (.A0(_3135_),
    .A1(\mem[27][21] ),
    .S(_4196_),
    .X(_4198_));
 sky130_fd_sc_hd__clkbuf_1 _8473_ (.A(_4198_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _8474_ (.A0(_3137_),
    .A1(\mem[27][22] ),
    .S(_4196_),
    .X(_4199_));
 sky130_fd_sc_hd__clkbuf_1 _8475_ (.A(_4199_),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _8476_ (.A0(_3139_),
    .A1(\mem[27][23] ),
    .S(_4196_),
    .X(_4200_));
 sky130_fd_sc_hd__clkbuf_1 _8477_ (.A(_4200_),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _8478_ (.A0(_3141_),
    .A1(\mem[27][24] ),
    .S(_4196_),
    .X(_4201_));
 sky130_fd_sc_hd__clkbuf_1 _8479_ (.A(_4201_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _8480_ (.A0(_3143_),
    .A1(\mem[27][25] ),
    .S(_4196_),
    .X(_4202_));
 sky130_fd_sc_hd__clkbuf_1 _8481_ (.A(_4202_),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _8482_ (.A0(_3145_),
    .A1(\mem[27][26] ),
    .S(_4196_),
    .X(_4203_));
 sky130_fd_sc_hd__clkbuf_1 _8483_ (.A(_4203_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _8484_ (.A0(_3147_),
    .A1(\mem[27][27] ),
    .S(_4196_),
    .X(_4204_));
 sky130_fd_sc_hd__clkbuf_1 _8485_ (.A(_4204_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _8486_ (.A0(_3149_),
    .A1(\mem[27][28] ),
    .S(_4196_),
    .X(_4205_));
 sky130_fd_sc_hd__clkbuf_1 _8487_ (.A(_4205_),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _8488_ (.A0(_3151_),
    .A1(\mem[27][29] ),
    .S(_4196_),
    .X(_4206_));
 sky130_fd_sc_hd__clkbuf_1 _8489_ (.A(_4206_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _8490_ (.A0(_3153_),
    .A1(\mem[27][30] ),
    .S(_4173_),
    .X(_4207_));
 sky130_fd_sc_hd__clkbuf_1 _8491_ (.A(_4207_),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _8492_ (.A0(_3155_),
    .A1(\mem[27][31] ),
    .S(_4173_),
    .X(_4208_));
 sky130_fd_sc_hd__clkbuf_1 _8493_ (.A(_4208_),
    .X(_0895_));
 sky130_fd_sc_hd__and3_4 _8494_ (.A(_3745_),
    .B(_3598_),
    .C(_3302_),
    .X(_4209_));
 sky130_fd_sc_hd__buf_6 _8495_ (.A(_4209_),
    .X(_4210_));
 sky130_fd_sc_hd__mux2_1 _8496_ (.A0(\mem[28][0] ),
    .A1(net18),
    .S(_4210_),
    .X(_4211_));
 sky130_fd_sc_hd__clkbuf_1 _8497_ (.A(_4211_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _8498_ (.A0(\mem[28][1] ),
    .A1(net29),
    .S(_4210_),
    .X(_4212_));
 sky130_fd_sc_hd__clkbuf_1 _8499_ (.A(_4212_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _8500_ (.A0(\mem[28][2] ),
    .A1(net40),
    .S(_4210_),
    .X(_4213_));
 sky130_fd_sc_hd__clkbuf_1 _8501_ (.A(_4213_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _8502_ (.A0(\mem[28][3] ),
    .A1(net43),
    .S(_4210_),
    .X(_4214_));
 sky130_fd_sc_hd__clkbuf_1 _8503_ (.A(_4214_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _8504_ (.A0(\mem[28][4] ),
    .A1(net44),
    .S(_4210_),
    .X(_4215_));
 sky130_fd_sc_hd__clkbuf_1 _8505_ (.A(_4215_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _8506_ (.A0(\mem[28][5] ),
    .A1(net45),
    .S(_4210_),
    .X(_4216_));
 sky130_fd_sc_hd__clkbuf_1 _8507_ (.A(_4216_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _8508_ (.A0(\mem[28][6] ),
    .A1(net46),
    .S(_4210_),
    .X(_4217_));
 sky130_fd_sc_hd__clkbuf_1 _8509_ (.A(_4217_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _8510_ (.A0(\mem[28][7] ),
    .A1(net47),
    .S(_4210_),
    .X(_4218_));
 sky130_fd_sc_hd__clkbuf_1 _8511_ (.A(_4218_),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _8512_ (.A0(\mem[28][8] ),
    .A1(net48),
    .S(_4210_),
    .X(_4219_));
 sky130_fd_sc_hd__clkbuf_1 _8513_ (.A(_4219_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _8514_ (.A0(\mem[28][9] ),
    .A1(net49),
    .S(_4210_),
    .X(_4220_));
 sky130_fd_sc_hd__clkbuf_1 _8515_ (.A(_4220_),
    .X(_0905_));
 sky130_fd_sc_hd__buf_6 _8516_ (.A(_4209_),
    .X(_4221_));
 sky130_fd_sc_hd__mux2_1 _8517_ (.A0(\mem[28][10] ),
    .A1(net19),
    .S(_4221_),
    .X(_4222_));
 sky130_fd_sc_hd__clkbuf_1 _8518_ (.A(_4222_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _8519_ (.A0(\mem[28][11] ),
    .A1(net20),
    .S(_4221_),
    .X(_4223_));
 sky130_fd_sc_hd__clkbuf_1 _8520_ (.A(_4223_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _8521_ (.A0(\mem[28][12] ),
    .A1(net21),
    .S(_4221_),
    .X(_4224_));
 sky130_fd_sc_hd__clkbuf_1 _8522_ (.A(_4224_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _8523_ (.A0(\mem[28][13] ),
    .A1(net22),
    .S(_4221_),
    .X(_4225_));
 sky130_fd_sc_hd__clkbuf_1 _8524_ (.A(_4225_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _8525_ (.A0(\mem[28][14] ),
    .A1(net23),
    .S(_4221_),
    .X(_4226_));
 sky130_fd_sc_hd__clkbuf_1 _8526_ (.A(_4226_),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _8527_ (.A0(\mem[28][15] ),
    .A1(net24),
    .S(_4221_),
    .X(_4227_));
 sky130_fd_sc_hd__clkbuf_1 _8528_ (.A(_4227_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _8529_ (.A0(\mem[28][16] ),
    .A1(net25),
    .S(_4221_),
    .X(_4228_));
 sky130_fd_sc_hd__clkbuf_1 _8530_ (.A(_4228_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _8531_ (.A0(\mem[28][17] ),
    .A1(net26),
    .S(_4221_),
    .X(_4229_));
 sky130_fd_sc_hd__clkbuf_1 _8532_ (.A(_4229_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _8533_ (.A0(\mem[28][18] ),
    .A1(net27),
    .S(_4221_),
    .X(_4230_));
 sky130_fd_sc_hd__clkbuf_1 _8534_ (.A(_4230_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _8535_ (.A0(\mem[28][19] ),
    .A1(net28),
    .S(_4221_),
    .X(_4231_));
 sky130_fd_sc_hd__clkbuf_1 _8536_ (.A(_4231_),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_8 _8537_ (.A(_4209_),
    .X(_4232_));
 sky130_fd_sc_hd__mux2_1 _8538_ (.A0(\mem[28][20] ),
    .A1(net30),
    .S(_4232_),
    .X(_4233_));
 sky130_fd_sc_hd__clkbuf_1 _8539_ (.A(_4233_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _8540_ (.A0(\mem[28][21] ),
    .A1(net31),
    .S(_4232_),
    .X(_4234_));
 sky130_fd_sc_hd__clkbuf_1 _8541_ (.A(_4234_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _8542_ (.A0(\mem[28][22] ),
    .A1(net32),
    .S(_4232_),
    .X(_4235_));
 sky130_fd_sc_hd__clkbuf_1 _8543_ (.A(_4235_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _8544_ (.A0(\mem[28][23] ),
    .A1(net33),
    .S(_4232_),
    .X(_4236_));
 sky130_fd_sc_hd__clkbuf_1 _8545_ (.A(_4236_),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_1 _8546_ (.A0(\mem[28][24] ),
    .A1(net34),
    .S(_4232_),
    .X(_4237_));
 sky130_fd_sc_hd__clkbuf_1 _8547_ (.A(_4237_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _8548_ (.A0(\mem[28][25] ),
    .A1(net35),
    .S(_4232_),
    .X(_4238_));
 sky130_fd_sc_hd__clkbuf_1 _8549_ (.A(_4238_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _8550_ (.A0(\mem[28][26] ),
    .A1(net36),
    .S(_4232_),
    .X(_4239_));
 sky130_fd_sc_hd__clkbuf_1 _8551_ (.A(_4239_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _8552_ (.A0(\mem[28][27] ),
    .A1(net37),
    .S(_4232_),
    .X(_4240_));
 sky130_fd_sc_hd__clkbuf_1 _8553_ (.A(_4240_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _8554_ (.A0(\mem[28][28] ),
    .A1(net38),
    .S(_4232_),
    .X(_4241_));
 sky130_fd_sc_hd__clkbuf_1 _8555_ (.A(_4241_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _8556_ (.A0(\mem[28][29] ),
    .A1(net39),
    .S(_4232_),
    .X(_4242_));
 sky130_fd_sc_hd__clkbuf_1 _8557_ (.A(_4242_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _8558_ (.A0(\mem[28][30] ),
    .A1(net41),
    .S(_4209_),
    .X(_4243_));
 sky130_fd_sc_hd__clkbuf_1 _8559_ (.A(_4243_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _8560_ (.A0(\mem[28][31] ),
    .A1(net42),
    .S(_4209_),
    .X(_4244_));
 sky130_fd_sc_hd__clkbuf_1 _8561_ (.A(_4244_),
    .X(_0927_));
 sky130_fd_sc_hd__or3_4 _8562_ (.A(_3087_),
    .B(_3089_),
    .C(_3340_),
    .X(_4245_));
 sky130_fd_sc_hd__buf_6 _8563_ (.A(_4245_),
    .X(_4246_));
 sky130_fd_sc_hd__mux2_1 _8564_ (.A0(_3157_),
    .A1(\mem[29][0] ),
    .S(_4246_),
    .X(_4247_));
 sky130_fd_sc_hd__clkbuf_1 _8565_ (.A(_4247_),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _8566_ (.A0(_3164_),
    .A1(\mem[29][1] ),
    .S(_4246_),
    .X(_4248_));
 sky130_fd_sc_hd__clkbuf_1 _8567_ (.A(_4248_),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_1 _8568_ (.A0(_3166_),
    .A1(\mem[29][2] ),
    .S(_4246_),
    .X(_4249_));
 sky130_fd_sc_hd__clkbuf_1 _8569_ (.A(_4249_),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _8570_ (.A0(_3168_),
    .A1(\mem[29][3] ),
    .S(_4246_),
    .X(_4250_));
 sky130_fd_sc_hd__clkbuf_1 _8571_ (.A(_4250_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _8572_ (.A0(_3170_),
    .A1(\mem[29][4] ),
    .S(_4246_),
    .X(_4251_));
 sky130_fd_sc_hd__clkbuf_1 _8573_ (.A(_4251_),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _8574_ (.A0(_3172_),
    .A1(\mem[29][5] ),
    .S(_4246_),
    .X(_4252_));
 sky130_fd_sc_hd__clkbuf_1 _8575_ (.A(_4252_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _8576_ (.A0(_3174_),
    .A1(\mem[29][6] ),
    .S(_4246_),
    .X(_4253_));
 sky130_fd_sc_hd__clkbuf_1 _8577_ (.A(_4253_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _8578_ (.A0(_3176_),
    .A1(\mem[29][7] ),
    .S(_4246_),
    .X(_4254_));
 sky130_fd_sc_hd__clkbuf_1 _8579_ (.A(_4254_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _8580_ (.A0(_3178_),
    .A1(\mem[29][8] ),
    .S(_4246_),
    .X(_4255_));
 sky130_fd_sc_hd__clkbuf_1 _8581_ (.A(_4255_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _8582_ (.A0(_3180_),
    .A1(\mem[29][9] ),
    .S(_4246_),
    .X(_4256_));
 sky130_fd_sc_hd__clkbuf_1 _8583_ (.A(_4256_),
    .X(_0937_));
 sky130_fd_sc_hd__buf_6 _8584_ (.A(_4245_),
    .X(_4257_));
 sky130_fd_sc_hd__mux2_1 _8585_ (.A0(_3182_),
    .A1(\mem[29][10] ),
    .S(_4257_),
    .X(_4258_));
 sky130_fd_sc_hd__clkbuf_1 _8586_ (.A(_4258_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _8587_ (.A0(_3185_),
    .A1(\mem[29][11] ),
    .S(_4257_),
    .X(_4259_));
 sky130_fd_sc_hd__clkbuf_1 _8588_ (.A(_4259_),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _8589_ (.A0(_3187_),
    .A1(\mem[29][12] ),
    .S(_4257_),
    .X(_4260_));
 sky130_fd_sc_hd__clkbuf_1 _8590_ (.A(_4260_),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_1 _8591_ (.A0(_3189_),
    .A1(\mem[29][13] ),
    .S(_4257_),
    .X(_4261_));
 sky130_fd_sc_hd__clkbuf_1 _8592_ (.A(_4261_),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _8593_ (.A0(_3191_),
    .A1(\mem[29][14] ),
    .S(_4257_),
    .X(_4262_));
 sky130_fd_sc_hd__clkbuf_1 _8594_ (.A(_4262_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _8595_ (.A0(_3193_),
    .A1(\mem[29][15] ),
    .S(_4257_),
    .X(_4263_));
 sky130_fd_sc_hd__clkbuf_1 _8596_ (.A(_4263_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _8597_ (.A0(_3195_),
    .A1(\mem[29][16] ),
    .S(_4257_),
    .X(_4264_));
 sky130_fd_sc_hd__clkbuf_1 _8598_ (.A(_4264_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _8599_ (.A0(_3197_),
    .A1(\mem[29][17] ),
    .S(_4257_),
    .X(_4265_));
 sky130_fd_sc_hd__clkbuf_1 _8600_ (.A(_4265_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _8601_ (.A0(_3199_),
    .A1(\mem[29][18] ),
    .S(_4257_),
    .X(_4266_));
 sky130_fd_sc_hd__clkbuf_1 _8602_ (.A(_4266_),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_1 _8603_ (.A0(_3201_),
    .A1(\mem[29][19] ),
    .S(_4257_),
    .X(_4267_));
 sky130_fd_sc_hd__clkbuf_1 _8604_ (.A(_4267_),
    .X(_0947_));
 sky130_fd_sc_hd__buf_4 _8605_ (.A(_4245_),
    .X(_4268_));
 sky130_fd_sc_hd__mux2_1 _8606_ (.A0(_3203_),
    .A1(\mem[29][20] ),
    .S(_4268_),
    .X(_4269_));
 sky130_fd_sc_hd__clkbuf_1 _8607_ (.A(_4269_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _8608_ (.A0(_3206_),
    .A1(\mem[29][21] ),
    .S(_4268_),
    .X(_4270_));
 sky130_fd_sc_hd__clkbuf_1 _8609_ (.A(_4270_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _8610_ (.A0(_3208_),
    .A1(\mem[29][22] ),
    .S(_4268_),
    .X(_4271_));
 sky130_fd_sc_hd__clkbuf_1 _8611_ (.A(_4271_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _8612_ (.A0(_3210_),
    .A1(\mem[29][23] ),
    .S(_4268_),
    .X(_4272_));
 sky130_fd_sc_hd__clkbuf_1 _8613_ (.A(_4272_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _8614_ (.A0(_3212_),
    .A1(\mem[29][24] ),
    .S(_4268_),
    .X(_4273_));
 sky130_fd_sc_hd__clkbuf_1 _8615_ (.A(_4273_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _8616_ (.A0(_3214_),
    .A1(\mem[29][25] ),
    .S(_4268_),
    .X(_4274_));
 sky130_fd_sc_hd__clkbuf_1 _8617_ (.A(_4274_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _8618_ (.A0(_3216_),
    .A1(\mem[29][26] ),
    .S(_4268_),
    .X(_4275_));
 sky130_fd_sc_hd__clkbuf_1 _8619_ (.A(_4275_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _8620_ (.A0(_3218_),
    .A1(\mem[29][27] ),
    .S(_4268_),
    .X(_4276_));
 sky130_fd_sc_hd__clkbuf_1 _8621_ (.A(_4276_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _8622_ (.A0(_3220_),
    .A1(\mem[29][28] ),
    .S(_4268_),
    .X(_4277_));
 sky130_fd_sc_hd__clkbuf_1 _8623_ (.A(_4277_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _8624_ (.A0(_3222_),
    .A1(\mem[29][29] ),
    .S(_4268_),
    .X(_4278_));
 sky130_fd_sc_hd__clkbuf_1 _8625_ (.A(_4278_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _8626_ (.A0(_3224_),
    .A1(\mem[29][30] ),
    .S(_4245_),
    .X(_4279_));
 sky130_fd_sc_hd__clkbuf_1 _8627_ (.A(_4279_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _8628_ (.A0(_3226_),
    .A1(\mem[29][31] ),
    .S(_4245_),
    .X(_4280_));
 sky130_fd_sc_hd__clkbuf_1 _8629_ (.A(_4280_),
    .X(_0959_));
 sky130_fd_sc_hd__or3_4 _8630_ (.A(_3087_),
    .B(_3089_),
    .C(_3379_),
    .X(_4281_));
 sky130_fd_sc_hd__buf_6 _8631_ (.A(_4281_),
    .X(_4282_));
 sky130_fd_sc_hd__mux2_1 _8632_ (.A0(_3157_),
    .A1(\mem[30][0] ),
    .S(_4282_),
    .X(_4283_));
 sky130_fd_sc_hd__clkbuf_1 _8633_ (.A(_4283_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _8634_ (.A0(_3164_),
    .A1(\mem[30][1] ),
    .S(_4282_),
    .X(_4284_));
 sky130_fd_sc_hd__clkbuf_1 _8635_ (.A(_4284_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _8636_ (.A0(_3166_),
    .A1(\mem[30][2] ),
    .S(_4282_),
    .X(_4285_));
 sky130_fd_sc_hd__clkbuf_1 _8637_ (.A(_4285_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _8638_ (.A0(_3168_),
    .A1(\mem[30][3] ),
    .S(_4282_),
    .X(_4286_));
 sky130_fd_sc_hd__clkbuf_1 _8639_ (.A(_4286_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _8640_ (.A0(_3170_),
    .A1(\mem[30][4] ),
    .S(_4282_),
    .X(_4287_));
 sky130_fd_sc_hd__clkbuf_1 _8641_ (.A(_4287_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _8642_ (.A0(_3172_),
    .A1(\mem[30][5] ),
    .S(_4282_),
    .X(_4288_));
 sky130_fd_sc_hd__clkbuf_1 _8643_ (.A(_4288_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _8644_ (.A0(_3174_),
    .A1(\mem[30][6] ),
    .S(_4282_),
    .X(_4289_));
 sky130_fd_sc_hd__clkbuf_1 _8645_ (.A(_4289_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _8646_ (.A0(_3176_),
    .A1(\mem[30][7] ),
    .S(_4282_),
    .X(_4290_));
 sky130_fd_sc_hd__clkbuf_1 _8647_ (.A(_4290_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _8648_ (.A0(_3178_),
    .A1(\mem[30][8] ),
    .S(_4282_),
    .X(_4291_));
 sky130_fd_sc_hd__clkbuf_1 _8649_ (.A(_4291_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _8650_ (.A0(_3180_),
    .A1(\mem[30][9] ),
    .S(_4282_),
    .X(_4292_));
 sky130_fd_sc_hd__clkbuf_1 _8651_ (.A(_4292_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_8 _8652_ (.A(_4281_),
    .X(_4293_));
 sky130_fd_sc_hd__mux2_1 _8653_ (.A0(_3182_),
    .A1(\mem[30][10] ),
    .S(_4293_),
    .X(_4294_));
 sky130_fd_sc_hd__clkbuf_1 _8654_ (.A(_4294_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _8655_ (.A0(_3185_),
    .A1(\mem[30][11] ),
    .S(_4293_),
    .X(_4295_));
 sky130_fd_sc_hd__clkbuf_1 _8656_ (.A(_4295_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _8657_ (.A0(_3187_),
    .A1(\mem[30][12] ),
    .S(_4293_),
    .X(_4296_));
 sky130_fd_sc_hd__clkbuf_1 _8658_ (.A(_4296_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _8659_ (.A0(_3189_),
    .A1(\mem[30][13] ),
    .S(_4293_),
    .X(_4297_));
 sky130_fd_sc_hd__clkbuf_1 _8660_ (.A(_4297_),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _8661_ (.A0(_3191_),
    .A1(\mem[30][14] ),
    .S(_4293_),
    .X(_4298_));
 sky130_fd_sc_hd__clkbuf_1 _8662_ (.A(_4298_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _8663_ (.A0(_3193_),
    .A1(\mem[30][15] ),
    .S(_4293_),
    .X(_4299_));
 sky130_fd_sc_hd__clkbuf_1 _8664_ (.A(_4299_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _8665_ (.A0(_3195_),
    .A1(\mem[30][16] ),
    .S(_4293_),
    .X(_4300_));
 sky130_fd_sc_hd__clkbuf_1 _8666_ (.A(_4300_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _8667_ (.A0(_3197_),
    .A1(\mem[30][17] ),
    .S(_4293_),
    .X(_4301_));
 sky130_fd_sc_hd__clkbuf_1 _8668_ (.A(_4301_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _8669_ (.A0(_3199_),
    .A1(\mem[30][18] ),
    .S(_4293_),
    .X(_4302_));
 sky130_fd_sc_hd__clkbuf_1 _8670_ (.A(_4302_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _8671_ (.A0(_3201_),
    .A1(\mem[30][19] ),
    .S(_4293_),
    .X(_4303_));
 sky130_fd_sc_hd__clkbuf_1 _8672_ (.A(_4303_),
    .X(_0979_));
 sky130_fd_sc_hd__buf_4 _8673_ (.A(_4281_),
    .X(_4304_));
 sky130_fd_sc_hd__mux2_1 _8674_ (.A0(_3203_),
    .A1(\mem[30][20] ),
    .S(_4304_),
    .X(_4305_));
 sky130_fd_sc_hd__clkbuf_1 _8675_ (.A(_4305_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _8676_ (.A0(_3206_),
    .A1(\mem[30][21] ),
    .S(_4304_),
    .X(_4306_));
 sky130_fd_sc_hd__clkbuf_1 _8677_ (.A(_4306_),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _8678_ (.A0(_3208_),
    .A1(\mem[30][22] ),
    .S(_4304_),
    .X(_4307_));
 sky130_fd_sc_hd__clkbuf_1 _8679_ (.A(_4307_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _8680_ (.A0(_3210_),
    .A1(\mem[30][23] ),
    .S(_4304_),
    .X(_4308_));
 sky130_fd_sc_hd__clkbuf_1 _8681_ (.A(_4308_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _8682_ (.A0(_3212_),
    .A1(\mem[30][24] ),
    .S(_4304_),
    .X(_4309_));
 sky130_fd_sc_hd__clkbuf_1 _8683_ (.A(_4309_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _8684_ (.A0(_3214_),
    .A1(\mem[30][25] ),
    .S(_4304_),
    .X(_4310_));
 sky130_fd_sc_hd__clkbuf_1 _8685_ (.A(_4310_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _8686_ (.A0(_3216_),
    .A1(\mem[30][26] ),
    .S(_4304_),
    .X(_4311_));
 sky130_fd_sc_hd__clkbuf_1 _8687_ (.A(_4311_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _8688_ (.A0(_3218_),
    .A1(\mem[30][27] ),
    .S(_4304_),
    .X(_4312_));
 sky130_fd_sc_hd__clkbuf_1 _8689_ (.A(_4312_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _8690_ (.A0(_3220_),
    .A1(\mem[30][28] ),
    .S(_4304_),
    .X(_4313_));
 sky130_fd_sc_hd__clkbuf_1 _8691_ (.A(_4313_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _8692_ (.A0(_3222_),
    .A1(\mem[30][29] ),
    .S(_4304_),
    .X(_4314_));
 sky130_fd_sc_hd__clkbuf_1 _8693_ (.A(_4314_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _8694_ (.A0(_3224_),
    .A1(\mem[30][30] ),
    .S(_4281_),
    .X(_4315_));
 sky130_fd_sc_hd__clkbuf_1 _8695_ (.A(_4315_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _8696_ (.A0(_3226_),
    .A1(\mem[30][31] ),
    .S(_4281_),
    .X(_4316_));
 sky130_fd_sc_hd__clkbuf_1 _8697_ (.A(_4316_),
    .X(_0991_));
 sky130_fd_sc_hd__dfrtp_1 _8698_ (.CLK(clk),
    .D(_0000_),
    .RESET_B(net187),
    .Q(\mem[31][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8699_ (.CLK(clk),
    .D(_0001_),
    .RESET_B(net125),
    .Q(\mem[31][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8700_ (.CLK(clk),
    .D(_0002_),
    .RESET_B(net125),
    .Q(\mem[31][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8701_ (.CLK(clk),
    .D(_0003_),
    .RESET_B(net198),
    .Q(\mem[31][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8702_ (.CLK(clk),
    .D(_0004_),
    .RESET_B(net194),
    .Q(\mem[31][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8703_ (.CLK(clk),
    .D(_0005_),
    .RESET_B(net175),
    .Q(\mem[31][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8704_ (.CLK(clk),
    .D(_0006_),
    .RESET_B(net180),
    .Q(\mem[31][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8705_ (.CLK(clk),
    .D(_0007_),
    .RESET_B(net205),
    .Q(\mem[31][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8706_ (.CLK(clk),
    .D(_0008_),
    .RESET_B(net206),
    .Q(\mem[31][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8707_ (.CLK(clk),
    .D(_0009_),
    .RESET_B(net208),
    .Q(\mem[31][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8708_ (.CLK(clk),
    .D(_0010_),
    .RESET_B(net208),
    .Q(\mem[31][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8709_ (.CLK(clk),
    .D(_0011_),
    .RESET_B(net233),
    .Q(\mem[31][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8710_ (.CLK(clk),
    .D(_0012_),
    .RESET_B(net227),
    .Q(\mem[31][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8711_ (.CLK(clk),
    .D(_0013_),
    .RESET_B(net235),
    .Q(\mem[31][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8712_ (.CLK(clk),
    .D(_0014_),
    .RESET_B(net235),
    .Q(\mem[31][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8713_ (.CLK(clk),
    .D(_0015_),
    .RESET_B(net240),
    .Q(\mem[31][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8714_ (.CLK(clk),
    .D(_0016_),
    .RESET_B(net242),
    .Q(\mem[31][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8715_ (.CLK(clk),
    .D(_0017_),
    .RESET_B(net226),
    .Q(\mem[31][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8716_ (.CLK(clk),
    .D(_0018_),
    .RESET_B(net221),
    .Q(\mem[31][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8717_ (.CLK(clk),
    .D(_0019_),
    .RESET_B(net170),
    .Q(\mem[31][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8718_ (.CLK(clk),
    .D(_0020_),
    .RESET_B(net150),
    .Q(\mem[31][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8719_ (.CLK(clk),
    .D(_0021_),
    .RESET_B(net150),
    .Q(\mem[31][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8720_ (.CLK(clk),
    .D(_0022_),
    .RESET_B(net148),
    .Q(\mem[31][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8721_ (.CLK(clk),
    .D(_0023_),
    .RESET_B(net148),
    .Q(\mem[31][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8722_ (.CLK(clk),
    .D(_0024_),
    .RESET_B(net148),
    .Q(\mem[31][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8723_ (.CLK(clk),
    .D(_0025_),
    .RESET_B(net140),
    .Q(\mem[31][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8724_ (.CLK(clk),
    .D(_0026_),
    .RESET_B(net137),
    .Q(\mem[31][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8725_ (.CLK(clk),
    .D(_0027_),
    .RESET_B(net137),
    .Q(\mem[31][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8726_ (.CLK(clk),
    .D(_0028_),
    .RESET_B(net115),
    .Q(\mem[31][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8727_ (.CLK(clk),
    .D(_0029_),
    .RESET_B(net114),
    .Q(\mem[31][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8728_ (.CLK(clk),
    .D(_0030_),
    .RESET_B(net118),
    .Q(\mem[31][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8729_ (.CLK(clk),
    .D(_0031_),
    .RESET_B(net117),
    .Q(\mem[31][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8730_ (.CLK(clk),
    .D(_0032_),
    .RESET_B(net186),
    .Q(\mem[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8731_ (.CLK(clk),
    .D(_0033_),
    .RESET_B(net135),
    .Q(\mem[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8732_ (.CLK(clk),
    .D(_0034_),
    .RESET_B(net184),
    .Q(\mem[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8733_ (.CLK(clk),
    .D(_0035_),
    .RESET_B(net184),
    .Q(\mem[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8734_ (.CLK(clk),
    .D(_0036_),
    .RESET_B(net188),
    .Q(\mem[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8735_ (.CLK(clk),
    .D(_0037_),
    .RESET_B(net184),
    .Q(\mem[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8736_ (.CLK(clk),
    .D(_0038_),
    .RESET_B(net184),
    .Q(\mem[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8737_ (.CLK(clk),
    .D(_0039_),
    .RESET_B(net188),
    .Q(\mem[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8738_ (.CLK(clk),
    .D(_0040_),
    .RESET_B(net190),
    .Q(\mem[1][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8739_ (.CLK(clk),
    .D(_0041_),
    .RESET_B(net190),
    .Q(\mem[1][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8740_ (.CLK(clk),
    .D(_0042_),
    .RESET_B(net190),
    .Q(\mem[1][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8741_ (.CLK(clk),
    .D(_0043_),
    .RESET_B(net214),
    .Q(\mem[1][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8742_ (.CLK(clk),
    .D(_0044_),
    .RESET_B(net211),
    .Q(\mem[1][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8743_ (.CLK(clk),
    .D(_0045_),
    .RESET_B(net214),
    .Q(\mem[1][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8744_ (.CLK(clk),
    .D(_0046_),
    .RESET_B(net216),
    .Q(\mem[1][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8745_ (.CLK(clk),
    .D(_0047_),
    .RESET_B(net224),
    .Q(\mem[1][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8746_ (.CLK(clk),
    .D(_0048_),
    .RESET_B(net224),
    .Q(\mem[1][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8747_ (.CLK(clk),
    .D(_0049_),
    .RESET_B(net219),
    .Q(\mem[1][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8748_ (.CLK(clk),
    .D(_0050_),
    .RESET_B(net211),
    .Q(\mem[1][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8749_ (.CLK(clk),
    .D(_0051_),
    .RESET_B(net219),
    .Q(\mem[1][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8750_ (.CLK(clk),
    .D(_0052_),
    .RESET_B(net170),
    .Q(\mem[1][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8751_ (.CLK(clk),
    .D(_0053_),
    .RESET_B(net170),
    .Q(\mem[1][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8752_ (.CLK(clk),
    .D(_0054_),
    .RESET_B(net161),
    .Q(\mem[1][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8753_ (.CLK(clk),
    .D(_0055_),
    .RESET_B(net170),
    .Q(\mem[1][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8754_ (.CLK(clk),
    .D(_0056_),
    .RESET_B(net169),
    .Q(\mem[1][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8755_ (.CLK(clk),
    .D(_0057_),
    .RESET_B(net162),
    .Q(\mem[1][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8756_ (.CLK(clk),
    .D(_0058_),
    .RESET_B(net163),
    .Q(\mem[1][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8757_ (.CLK(clk),
    .D(_0059_),
    .RESET_B(net163),
    .Q(\mem[1][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8758_ (.CLK(clk),
    .D(_0060_),
    .RESET_B(net163),
    .Q(\mem[1][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8759_ (.CLK(clk),
    .D(_0061_),
    .RESET_B(net134),
    .Q(\mem[1][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8760_ (.CLK(clk),
    .D(_0062_),
    .RESET_B(net135),
    .Q(\mem[1][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8761_ (.CLK(clk),
    .D(_0063_),
    .RESET_B(net135),
    .Q(\mem[1][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8762_ (.CLK(clk),
    .D(_0064_),
    .RESET_B(net186),
    .Q(\mem[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8763_ (.CLK(clk),
    .D(_0065_),
    .RESET_B(net128),
    .Q(\mem[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8764_ (.CLK(clk),
    .D(_0066_),
    .RESET_B(net127),
    .Q(\mem[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8765_ (.CLK(clk),
    .D(_0067_),
    .RESET_B(net196),
    .Q(\mem[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8766_ (.CLK(clk),
    .D(_0068_),
    .RESET_B(net194),
    .Q(\mem[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8767_ (.CLK(clk),
    .D(_0069_),
    .RESET_B(net176),
    .Q(\mem[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8768_ (.CLK(clk),
    .D(_0070_),
    .RESET_B(net177),
    .Q(\mem[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8769_ (.CLK(clk),
    .D(_0071_),
    .RESET_B(net196),
    .Q(\mem[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8770_ (.CLK(clk),
    .D(_0072_),
    .RESET_B(net201),
    .Q(\mem[2][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8771_ (.CLK(clk),
    .D(_0073_),
    .RESET_B(net203),
    .Q(\mem[2][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8772_ (.CLK(clk),
    .D(_0074_),
    .RESET_B(net229),
    .Q(\mem[2][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8773_ (.CLK(clk),
    .D(_0075_),
    .RESET_B(net229),
    .Q(\mem[2][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8774_ (.CLK(clk),
    .D(_0076_),
    .RESET_B(net224),
    .Q(\mem[2][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8775_ (.CLK(clk),
    .D(_0077_),
    .RESET_B(net231),
    .Q(\mem[2][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8776_ (.CLK(clk),
    .D(_0078_),
    .RESET_B(net231),
    .Q(\mem[2][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8777_ (.CLK(clk),
    .D(_0079_),
    .RESET_B(net238),
    .Q(\mem[2][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8778_ (.CLK(clk),
    .D(_0080_),
    .RESET_B(net238),
    .Q(\mem[2][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8779_ (.CLK(clk),
    .D(_0081_),
    .RESET_B(net220),
    .Q(\mem[2][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8780_ (.CLK(clk),
    .D(_0082_),
    .RESET_B(net161),
    .Q(\mem[2][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8781_ (.CLK(clk),
    .D(_0083_),
    .RESET_B(net169),
    .Q(\mem[2][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8782_ (.CLK(clk),
    .D(_0084_),
    .RESET_B(net166),
    .Q(\mem[2][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8783_ (.CLK(clk),
    .D(_0085_),
    .RESET_B(net154),
    .Q(\mem[2][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8784_ (.CLK(clk),
    .D(_0086_),
    .RESET_B(net145),
    .Q(\mem[2][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8785_ (.CLK(clk),
    .D(_0087_),
    .RESET_B(net155),
    .Q(\mem[2][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8786_ (.CLK(clk),
    .D(_0088_),
    .RESET_B(net152),
    .Q(\mem[2][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8787_ (.CLK(clk),
    .D(_0089_),
    .RESET_B(net146),
    .Q(\mem[2][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8788_ (.CLK(clk),
    .D(_0090_),
    .RESET_B(net144),
    .Q(\mem[2][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8789_ (.CLK(clk),
    .D(_0091_),
    .RESET_B(net144),
    .Q(\mem[2][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8790_ (.CLK(clk),
    .D(_0092_),
    .RESET_B(net144),
    .Q(\mem[2][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8791_ (.CLK(clk),
    .D(_0093_),
    .RESET_B(net131),
    .Q(\mem[2][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8792_ (.CLK(clk),
    .D(_0094_),
    .RESET_B(net122),
    .Q(\mem[2][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8793_ (.CLK(clk),
    .D(_0095_),
    .RESET_B(net122),
    .Q(\mem[2][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8794_ (.CLK(clk),
    .D(_0096_),
    .RESET_B(net186),
    .Q(\mem[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8795_ (.CLK(clk),
    .D(_0097_),
    .RESET_B(net135),
    .Q(\mem[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8796_ (.CLK(clk),
    .D(_0098_),
    .RESET_B(net184),
    .Q(\mem[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8797_ (.CLK(clk),
    .D(_0099_),
    .RESET_B(net185),
    .Q(\mem[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8798_ (.CLK(clk),
    .D(_0100_),
    .RESET_B(net188),
    .Q(\mem[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8799_ (.CLK(clk),
    .D(_0101_),
    .RESET_B(net184),
    .Q(\mem[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8800_ (.CLK(clk),
    .D(_0102_),
    .RESET_B(net185),
    .Q(\mem[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8801_ (.CLK(clk),
    .D(_0103_),
    .RESET_B(net188),
    .Q(\mem[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8802_ (.CLK(clk),
    .D(_0104_),
    .RESET_B(net190),
    .Q(\mem[3][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8803_ (.CLK(clk),
    .D(_0105_),
    .RESET_B(net190),
    .Q(\mem[3][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8804_ (.CLK(clk),
    .D(_0106_),
    .RESET_B(net214),
    .Q(\mem[3][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8805_ (.CLK(clk),
    .D(_0107_),
    .RESET_B(net214),
    .Q(\mem[3][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8806_ (.CLK(clk),
    .D(_0108_),
    .RESET_B(net211),
    .Q(\mem[3][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8807_ (.CLK(clk),
    .D(_0109_),
    .RESET_B(net214),
    .Q(\mem[3][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8808_ (.CLK(clk),
    .D(_0110_),
    .RESET_B(net216),
    .Q(\mem[3][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8809_ (.CLK(clk),
    .D(_0111_),
    .RESET_B(net224),
    .Q(\mem[3][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8810_ (.CLK(clk),
    .D(_0112_),
    .RESET_B(net224),
    .Q(\mem[3][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8811_ (.CLK(clk),
    .D(_0113_),
    .RESET_B(net220),
    .Q(\mem[3][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8812_ (.CLK(clk),
    .D(_0114_),
    .RESET_B(net213),
    .Q(\mem[3][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8813_ (.CLK(clk),
    .D(_0115_),
    .RESET_B(net169),
    .Q(\mem[3][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8814_ (.CLK(clk),
    .D(_0116_),
    .RESET_B(net170),
    .Q(\mem[3][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8815_ (.CLK(clk),
    .D(_0117_),
    .RESET_B(net170),
    .Q(\mem[3][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8816_ (.CLK(clk),
    .D(_0118_),
    .RESET_B(net161),
    .Q(\mem[3][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8817_ (.CLK(clk),
    .D(_0119_),
    .RESET_B(net170),
    .Q(\mem[3][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8818_ (.CLK(clk),
    .D(_0120_),
    .RESET_B(net162),
    .Q(\mem[3][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8819_ (.CLK(clk),
    .D(_0121_),
    .RESET_B(net161),
    .Q(\mem[3][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8820_ (.CLK(clk),
    .D(_0122_),
    .RESET_B(net163),
    .Q(\mem[3][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8821_ (.CLK(clk),
    .D(_0123_),
    .RESET_B(net163),
    .Q(\mem[3][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8822_ (.CLK(clk),
    .D(_0124_),
    .RESET_B(net163),
    .Q(\mem[3][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8823_ (.CLK(clk),
    .D(_0125_),
    .RESET_B(net134),
    .Q(\mem[3][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8824_ (.CLK(clk),
    .D(_0126_),
    .RESET_B(net127),
    .Q(\mem[3][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8825_ (.CLK(clk),
    .D(_0127_),
    .RESET_B(net127),
    .Q(\mem[3][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8826_ (.CLK(clk),
    .D(_0128_),
    .RESET_B(net213),
    .Q(\mem[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8827_ (.CLK(clk),
    .D(_0129_),
    .RESET_B(net123),
    .Q(\mem[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8828_ (.CLK(clk),
    .D(_0130_),
    .RESET_B(net124),
    .Q(\mem[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8829_ (.CLK(clk),
    .D(_0131_),
    .RESET_B(net196),
    .Q(\mem[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8830_ (.CLK(clk),
    .D(_0132_),
    .RESET_B(net180),
    .Q(\mem[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8831_ (.CLK(clk),
    .D(_0133_),
    .RESET_B(net177),
    .Q(\mem[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8832_ (.CLK(clk),
    .D(_0134_),
    .RESET_B(net179),
    .Q(\mem[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8833_ (.CLK(clk),
    .D(_0135_),
    .RESET_B(net201),
    .Q(\mem[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8834_ (.CLK(clk),
    .D(_0136_),
    .RESET_B(net201),
    .Q(\mem[4][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8835_ (.CLK(clk),
    .D(_0137_),
    .RESET_B(net203),
    .Q(\mem[4][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8836_ (.CLK(clk),
    .D(_0138_),
    .RESET_B(net203),
    .Q(\mem[4][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8837_ (.CLK(clk),
    .D(_0139_),
    .RESET_B(net229),
    .Q(\mem[4][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8838_ (.CLK(clk),
    .D(_0140_),
    .RESET_B(net226),
    .Q(\mem[4][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8839_ (.CLK(clk),
    .D(_0141_),
    .RESET_B(net229),
    .Q(\mem[4][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8840_ (.CLK(clk),
    .D(_0142_),
    .RESET_B(net231),
    .Q(\mem[4][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8841_ (.CLK(clk),
    .D(_0143_),
    .RESET_B(net240),
    .Q(\mem[4][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8842_ (.CLK(clk),
    .D(_0144_),
    .RESET_B(net238),
    .Q(\mem[4][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8843_ (.CLK(clk),
    .D(_0145_),
    .RESET_B(net221),
    .Q(\mem[4][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8844_ (.CLK(clk),
    .D(_0146_),
    .RESET_B(net161),
    .Q(\mem[4][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8845_ (.CLK(clk),
    .D(_0147_),
    .RESET_B(net221),
    .Q(\mem[4][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8846_ (.CLK(clk),
    .D(_0148_),
    .RESET_B(net166),
    .Q(\mem[4][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8847_ (.CLK(clk),
    .D(_0149_),
    .RESET_B(net152),
    .Q(\mem[4][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8848_ (.CLK(clk),
    .D(_0150_),
    .RESET_B(net145),
    .Q(\mem[4][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8849_ (.CLK(clk),
    .D(_0151_),
    .RESET_B(net153),
    .Q(\mem[4][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8850_ (.CLK(clk),
    .D(_0152_),
    .RESET_B(net152),
    .Q(\mem[4][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8851_ (.CLK(clk),
    .D(_0153_),
    .RESET_B(net145),
    .Q(\mem[4][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8852_ (.CLK(clk),
    .D(_0154_),
    .RESET_B(net143),
    .Q(\mem[4][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8853_ (.CLK(clk),
    .D(_0155_),
    .RESET_B(net143),
    .Q(\mem[4][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8854_ (.CLK(clk),
    .D(_0156_),
    .RESET_B(net118),
    .Q(\mem[4][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8855_ (.CLK(clk),
    .D(_0157_),
    .RESET_B(net131),
    .Q(\mem[4][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8856_ (.CLK(clk),
    .D(_0158_),
    .RESET_B(net122),
    .Q(\mem[4][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8857_ (.CLK(clk),
    .D(_0159_),
    .RESET_B(net122),
    .Q(\mem[4][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8858_ (.CLK(clk),
    .D(_0160_),
    .RESET_B(net187),
    .Q(\mem[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8859_ (.CLK(clk),
    .D(_0161_),
    .RESET_B(net135),
    .Q(\mem[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8860_ (.CLK(clk),
    .D(_0162_),
    .RESET_B(net184),
    .Q(\mem[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8861_ (.CLK(clk),
    .D(_0163_),
    .RESET_B(net185),
    .Q(\mem[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8862_ (.CLK(clk),
    .D(_0164_),
    .RESET_B(net188),
    .Q(\mem[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8863_ (.CLK(clk),
    .D(_0165_),
    .RESET_B(net185),
    .Q(\mem[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8864_ (.CLK(clk),
    .D(_0166_),
    .RESET_B(net185),
    .Q(\mem[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8865_ (.CLK(clk),
    .D(_0167_),
    .RESET_B(net188),
    .Q(\mem[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8866_ (.CLK(clk),
    .D(_0168_),
    .RESET_B(net188),
    .Q(\mem[5][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8867_ (.CLK(clk),
    .D(_0169_),
    .RESET_B(net190),
    .Q(\mem[5][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8868_ (.CLK(clk),
    .D(_0170_),
    .RESET_B(net190),
    .Q(\mem[5][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8869_ (.CLK(clk),
    .D(_0171_),
    .RESET_B(net214),
    .Q(\mem[5][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8870_ (.CLK(clk),
    .D(_0172_),
    .RESET_B(net213),
    .Q(\mem[5][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8871_ (.CLK(clk),
    .D(_0173_),
    .RESET_B(net214),
    .Q(\mem[5][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8872_ (.CLK(clk),
    .D(_0174_),
    .RESET_B(net216),
    .Q(\mem[5][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8873_ (.CLK(clk),
    .D(_0175_),
    .RESET_B(net224),
    .Q(\mem[5][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8874_ (.CLK(clk),
    .D(_0176_),
    .RESET_B(net224),
    .Q(\mem[5][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8875_ (.CLK(clk),
    .D(_0177_),
    .RESET_B(net220),
    .Q(\mem[5][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8876_ (.CLK(clk),
    .D(_0178_),
    .RESET_B(net213),
    .Q(\mem[5][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8877_ (.CLK(clk),
    .D(_0179_),
    .RESET_B(net219),
    .Q(\mem[5][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8878_ (.CLK(clk),
    .D(_0180_),
    .RESET_B(net170),
    .Q(\mem[5][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8879_ (.CLK(clk),
    .D(_0181_),
    .RESET_B(net170),
    .Q(\mem[5][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8880_ (.CLK(clk),
    .D(_0182_),
    .RESET_B(net162),
    .Q(\mem[5][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8881_ (.CLK(clk),
    .D(_0183_),
    .RESET_B(net170),
    .Q(\mem[5][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8882_ (.CLK(clk),
    .D(_0184_),
    .RESET_B(net169),
    .Q(\mem[5][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8883_ (.CLK(clk),
    .D(_0185_),
    .RESET_B(net162),
    .Q(\mem[5][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8884_ (.CLK(clk),
    .D(_0186_),
    .RESET_B(net163),
    .Q(\mem[5][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8885_ (.CLK(clk),
    .D(_0187_),
    .RESET_B(net163),
    .Q(\mem[5][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8886_ (.CLK(clk),
    .D(_0188_),
    .RESET_B(net134),
    .Q(\mem[5][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8887_ (.CLK(clk),
    .D(_0189_),
    .RESET_B(net134),
    .Q(\mem[5][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8888_ (.CLK(clk),
    .D(_0190_),
    .RESET_B(net134),
    .Q(\mem[5][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8889_ (.CLK(clk),
    .D(_0191_),
    .RESET_B(net135),
    .Q(\mem[5][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8890_ (.CLK(clk),
    .D(_0192_),
    .RESET_B(net187),
    .Q(\mem[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8891_ (.CLK(clk),
    .D(_0193_),
    .RESET_B(net176),
    .Q(\mem[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8892_ (.CLK(clk),
    .D(_0194_),
    .RESET_B(net174),
    .Q(\mem[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8893_ (.CLK(clk),
    .D(_0195_),
    .RESET_B(net197),
    .Q(\mem[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8894_ (.CLK(clk),
    .D(_0196_),
    .RESET_B(net180),
    .Q(\mem[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8895_ (.CLK(clk),
    .D(_0197_),
    .RESET_B(net174),
    .Q(\mem[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8896_ (.CLK(clk),
    .D(_0198_),
    .RESET_B(net179),
    .Q(\mem[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8897_ (.CLK(clk),
    .D(_0199_),
    .RESET_B(net197),
    .Q(\mem[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8898_ (.CLK(clk),
    .D(_0200_),
    .RESET_B(net202),
    .Q(\mem[6][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8899_ (.CLK(clk),
    .D(_0201_),
    .RESET_B(net203),
    .Q(\mem[6][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8900_ (.CLK(clk),
    .D(_0202_),
    .RESET_B(net204),
    .Q(\mem[6][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8901_ (.CLK(clk),
    .D(_0203_),
    .RESET_B(net234),
    .Q(\mem[6][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8902_ (.CLK(clk),
    .D(_0204_),
    .RESET_B(net226),
    .Q(\mem[6][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8903_ (.CLK(clk),
    .D(_0205_),
    .RESET_B(net234),
    .Q(\mem[6][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8904_ (.CLK(clk),
    .D(_0206_),
    .RESET_B(net236),
    .Q(\mem[6][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8905_ (.CLK(clk),
    .D(_0207_),
    .RESET_B(net240),
    .Q(\mem[6][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8906_ (.CLK(clk),
    .D(_0208_),
    .RESET_B(net242),
    .Q(\mem[6][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8907_ (.CLK(clk),
    .D(_0209_),
    .RESET_B(net222),
    .Q(\mem[6][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8908_ (.CLK(clk),
    .D(_0210_),
    .RESET_B(net211),
    .Q(\mem[6][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8909_ (.CLK(clk),
    .D(_0211_),
    .RESET_B(net221),
    .Q(\mem[6][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8910_ (.CLK(clk),
    .D(_0212_),
    .RESET_B(net166),
    .Q(\mem[6][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8911_ (.CLK(clk),
    .D(_0213_),
    .RESET_B(net154),
    .Q(\mem[6][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8912_ (.CLK(clk),
    .D(_0214_),
    .RESET_B(net145),
    .Q(\mem[6][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8913_ (.CLK(clk),
    .D(_0215_),
    .RESET_B(net155),
    .Q(\mem[6][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8914_ (.CLK(clk),
    .D(_0216_),
    .RESET_B(net152),
    .Q(\mem[6][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8915_ (.CLK(clk),
    .D(_0217_),
    .RESET_B(net145),
    .Q(\mem[6][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8916_ (.CLK(clk),
    .D(_0218_),
    .RESET_B(net143),
    .Q(\mem[6][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8917_ (.CLK(clk),
    .D(_0219_),
    .RESET_B(net143),
    .Q(\mem[6][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8918_ (.CLK(clk),
    .D(_0220_),
    .RESET_B(net118),
    .Q(\mem[6][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8919_ (.CLK(clk),
    .D(_0221_),
    .RESET_B(net119),
    .Q(\mem[6][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8920_ (.CLK(clk),
    .D(_0222_),
    .RESET_B(net130),
    .Q(\mem[6][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8921_ (.CLK(clk),
    .D(_0223_),
    .RESET_B(net130),
    .Q(\mem[6][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8922_ (.CLK(clk),
    .D(_0224_),
    .RESET_B(net187),
    .Q(\mem[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8923_ (.CLK(clk),
    .D(_0225_),
    .RESET_B(net126),
    .Q(\mem[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8924_ (.CLK(clk),
    .D(_0226_),
    .RESET_B(net174),
    .Q(\mem[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8925_ (.CLK(clk),
    .D(_0227_),
    .RESET_B(net199),
    .Q(\mem[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8926_ (.CLK(clk),
    .D(_0228_),
    .RESET_B(net194),
    .Q(\mem[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8927_ (.CLK(clk),
    .D(_0229_),
    .RESET_B(net174),
    .Q(\mem[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8928_ (.CLK(clk),
    .D(_0230_),
    .RESET_B(net179),
    .Q(\mem[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8929_ (.CLK(clk),
    .D(_0231_),
    .RESET_B(net206),
    .Q(\mem[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8930_ (.CLK(clk),
    .D(_0232_),
    .RESET_B(net206),
    .Q(\mem[7][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8931_ (.CLK(clk),
    .D(_0233_),
    .RESET_B(net208),
    .Q(\mem[7][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8932_ (.CLK(clk),
    .D(_0234_),
    .RESET_B(net208),
    .Q(\mem[7][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8933_ (.CLK(clk),
    .D(_0235_),
    .RESET_B(net233),
    .Q(\mem[7][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8934_ (.CLK(clk),
    .D(_0236_),
    .RESET_B(net227),
    .Q(\mem[7][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8935_ (.CLK(clk),
    .D(_0237_),
    .RESET_B(net233),
    .Q(\mem[7][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8936_ (.CLK(clk),
    .D(_0238_),
    .RESET_B(net235),
    .Q(\mem[7][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8937_ (.CLK(clk),
    .D(_0239_),
    .RESET_B(net240),
    .Q(\mem[7][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8938_ (.CLK(clk),
    .D(_0240_),
    .RESET_B(net243),
    .Q(\mem[7][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8939_ (.CLK(clk),
    .D(_0241_),
    .RESET_B(net222),
    .Q(\mem[7][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8940_ (.CLK(clk),
    .D(_0242_),
    .RESET_B(net221),
    .Q(\mem[7][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8941_ (.CLK(clk),
    .D(_0243_),
    .RESET_B(net221),
    .Q(\mem[7][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8942_ (.CLK(clk),
    .D(_0244_),
    .RESET_B(net154),
    .Q(\mem[7][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8943_ (.CLK(clk),
    .D(_0245_),
    .RESET_B(net149),
    .Q(\mem[7][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8944_ (.CLK(clk),
    .D(_0246_),
    .RESET_B(net140),
    .Q(\mem[7][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8945_ (.CLK(clk),
    .D(_0247_),
    .RESET_B(net150),
    .Q(\mem[7][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8946_ (.CLK(clk),
    .D(_0248_),
    .RESET_B(net148),
    .Q(\mem[7][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8947_ (.CLK(clk),
    .D(_0249_),
    .RESET_B(net140),
    .Q(\mem[7][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8948_ (.CLK(clk),
    .D(_0250_),
    .RESET_B(net137),
    .Q(\mem[7][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8949_ (.CLK(clk),
    .D(_0251_),
    .RESET_B(net137),
    .Q(\mem[7][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8950_ (.CLK(clk),
    .D(_0252_),
    .RESET_B(net115),
    .Q(\mem[7][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8951_ (.CLK(clk),
    .D(_0253_),
    .RESET_B(net114),
    .Q(\mem[7][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8952_ (.CLK(clk),
    .D(_0254_),
    .RESET_B(net117),
    .Q(\mem[7][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8953_ (.CLK(clk),
    .D(_0255_),
    .RESET_B(net117),
    .Q(\mem[7][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8954_ (.CLK(clk),
    .D(_0256_),
    .RESET_B(net186),
    .Q(\mem[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8955_ (.CLK(clk),
    .D(_0257_),
    .RESET_B(net176),
    .Q(\mem[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8956_ (.CLK(clk),
    .D(_0258_),
    .RESET_B(net176),
    .Q(\mem[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8957_ (.CLK(clk),
    .D(_0259_),
    .RESET_B(net197),
    .Q(\mem[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8958_ (.CLK(clk),
    .D(_0260_),
    .RESET_B(net194),
    .Q(\mem[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8959_ (.CLK(clk),
    .D(_0261_),
    .RESET_B(net175),
    .Q(\mem[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8960_ (.CLK(clk),
    .D(_0262_),
    .RESET_B(net179),
    .Q(\mem[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8961_ (.CLK(clk),
    .D(_0263_),
    .RESET_B(net197),
    .Q(\mem[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8962_ (.CLK(clk),
    .D(_0264_),
    .RESET_B(net202),
    .Q(\mem[8][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8963_ (.CLK(clk),
    .D(_0265_),
    .RESET_B(net204),
    .Q(\mem[8][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8964_ (.CLK(clk),
    .D(_0266_),
    .RESET_B(net204),
    .Q(\mem[8][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8965_ (.CLK(clk),
    .D(_0267_),
    .RESET_B(net229),
    .Q(\mem[8][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8966_ (.CLK(clk),
    .D(_0268_),
    .RESET_B(net226),
    .Q(\mem[8][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8967_ (.CLK(clk),
    .D(_0269_),
    .RESET_B(net234),
    .Q(\mem[8][13] ));
 sky130_fd_sc_hd__dfrtp_1 _8968_ (.CLK(clk),
    .D(_0270_),
    .RESET_B(net236),
    .Q(\mem[8][14] ));
 sky130_fd_sc_hd__dfrtp_1 _8969_ (.CLK(clk),
    .D(_0271_),
    .RESET_B(net240),
    .Q(\mem[8][15] ));
 sky130_fd_sc_hd__dfrtp_1 _8970_ (.CLK(clk),
    .D(_0272_),
    .RESET_B(net238),
    .Q(\mem[8][16] ));
 sky130_fd_sc_hd__dfrtp_1 _8971_ (.CLK(clk),
    .D(_0273_),
    .RESET_B(net222),
    .Q(\mem[8][17] ));
 sky130_fd_sc_hd__dfrtp_1 _8972_ (.CLK(clk),
    .D(_0274_),
    .RESET_B(net211),
    .Q(\mem[8][18] ));
 sky130_fd_sc_hd__dfrtp_1 _8973_ (.CLK(clk),
    .D(_0275_),
    .RESET_B(net221),
    .Q(\mem[8][19] ));
 sky130_fd_sc_hd__dfrtp_1 _8974_ (.CLK(clk),
    .D(_0276_),
    .RESET_B(net167),
    .Q(\mem[8][20] ));
 sky130_fd_sc_hd__dfrtp_1 _8975_ (.CLK(clk),
    .D(_0277_),
    .RESET_B(net154),
    .Q(\mem[8][21] ));
 sky130_fd_sc_hd__dfrtp_1 _8976_ (.CLK(clk),
    .D(_0278_),
    .RESET_B(net145),
    .Q(\mem[8][22] ));
 sky130_fd_sc_hd__dfrtp_1 _8977_ (.CLK(clk),
    .D(_0279_),
    .RESET_B(net155),
    .Q(\mem[8][23] ));
 sky130_fd_sc_hd__dfrtp_1 _8978_ (.CLK(clk),
    .D(_0280_),
    .RESET_B(net152),
    .Q(\mem[8][24] ));
 sky130_fd_sc_hd__dfrtp_1 _8979_ (.CLK(clk),
    .D(_0281_),
    .RESET_B(net145),
    .Q(\mem[8][25] ));
 sky130_fd_sc_hd__dfrtp_1 _8980_ (.CLK(clk),
    .D(_0282_),
    .RESET_B(net143),
    .Q(\mem[8][26] ));
 sky130_fd_sc_hd__dfrtp_1 _8981_ (.CLK(clk),
    .D(_0283_),
    .RESET_B(net143),
    .Q(\mem[8][27] ));
 sky130_fd_sc_hd__dfrtp_1 _8982_ (.CLK(clk),
    .D(_0284_),
    .RESET_B(net143),
    .Q(\mem[8][28] ));
 sky130_fd_sc_hd__dfrtp_1 _8983_ (.CLK(clk),
    .D(_0285_),
    .RESET_B(net131),
    .Q(\mem[8][29] ));
 sky130_fd_sc_hd__dfrtp_1 _8984_ (.CLK(clk),
    .D(_0286_),
    .RESET_B(net130),
    .Q(\mem[8][30] ));
 sky130_fd_sc_hd__dfrtp_1 _8985_ (.CLK(clk),
    .D(_0287_),
    .RESET_B(net130),
    .Q(\mem[8][31] ));
 sky130_fd_sc_hd__dfrtp_1 _8986_ (.CLK(clk),
    .D(_0288_),
    .RESET_B(net134),
    .Q(\mem[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8987_ (.CLK(clk),
    .D(_0289_),
    .RESET_B(net126),
    .Q(\mem[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8988_ (.CLK(clk),
    .D(_0290_),
    .RESET_B(net174),
    .Q(\mem[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _8989_ (.CLK(clk),
    .D(_0291_),
    .RESET_B(net199),
    .Q(\mem[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _8990_ (.CLK(clk),
    .D(_0292_),
    .RESET_B(net194),
    .Q(\mem[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _8991_ (.CLK(clk),
    .D(_0293_),
    .RESET_B(net175),
    .Q(\mem[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _8992_ (.CLK(clk),
    .D(_0294_),
    .RESET_B(net179),
    .Q(\mem[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _8993_ (.CLK(clk),
    .D(_0295_),
    .RESET_B(net206),
    .Q(\mem[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _8994_ (.CLK(clk),
    .D(_0296_),
    .RESET_B(net206),
    .Q(\mem[9][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8995_ (.CLK(clk),
    .D(_0297_),
    .RESET_B(net208),
    .Q(\mem[9][9] ));
 sky130_fd_sc_hd__dfrtp_1 _8996_ (.CLK(clk),
    .D(_0298_),
    .RESET_B(net208),
    .Q(\mem[9][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8997_ (.CLK(clk),
    .D(_0299_),
    .RESET_B(net233),
    .Q(\mem[9][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8998_ (.CLK(clk),
    .D(_0300_),
    .RESET_B(net227),
    .Q(\mem[9][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8999_ (.CLK(clk),
    .D(_0301_),
    .RESET_B(net233),
    .Q(\mem[9][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9000_ (.CLK(clk),
    .D(_0302_),
    .RESET_B(net235),
    .Q(\mem[9][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9001_ (.CLK(clk),
    .D(_0303_),
    .RESET_B(net241),
    .Q(\mem[9][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9002_ (.CLK(clk),
    .D(_0304_),
    .RESET_B(net243),
    .Q(\mem[9][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9003_ (.CLK(clk),
    .D(_0305_),
    .RESET_B(net222),
    .Q(\mem[9][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9004_ (.CLK(clk),
    .D(_0306_),
    .RESET_B(net222),
    .Q(\mem[9][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9005_ (.CLK(clk),
    .D(_0307_),
    .RESET_B(net171),
    .Q(\mem[9][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9006_ (.CLK(clk),
    .D(_0308_),
    .RESET_B(net150),
    .Q(\mem[9][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9007_ (.CLK(clk),
    .D(_0309_),
    .RESET_B(net150),
    .Q(\mem[9][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9008_ (.CLK(clk),
    .D(_0310_),
    .RESET_B(net140),
    .Q(\mem[9][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9009_ (.CLK(clk),
    .D(_0311_),
    .RESET_B(net150),
    .Q(\mem[9][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9010_ (.CLK(clk),
    .D(_0312_),
    .RESET_B(net148),
    .Q(\mem[9][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9011_ (.CLK(clk),
    .D(_0313_),
    .RESET_B(net140),
    .Q(\mem[9][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9012_ (.CLK(clk),
    .D(_0314_),
    .RESET_B(net137),
    .Q(\mem[9][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9013_ (.CLK(clk),
    .D(_0315_),
    .RESET_B(net137),
    .Q(\mem[9][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9014_ (.CLK(clk),
    .D(_0316_),
    .RESET_B(net115),
    .Q(\mem[9][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9015_ (.CLK(clk),
    .D(_0317_),
    .RESET_B(net114),
    .Q(\mem[9][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9016_ (.CLK(clk),
    .D(_0318_),
    .RESET_B(net117),
    .Q(\mem[9][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9017_ (.CLK(clk),
    .D(_0319_),
    .RESET_B(net117),
    .Q(\mem[9][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9018_ (.CLK(clk),
    .D(_0320_),
    .RESET_B(net134),
    .Q(\mem[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9019_ (.CLK(clk),
    .D(_0321_),
    .RESET_B(net128),
    .Q(\mem[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9020_ (.CLK(clk),
    .D(_0322_),
    .RESET_B(net127),
    .Q(\mem[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9021_ (.CLK(clk),
    .D(_0323_),
    .RESET_B(net196),
    .Q(\mem[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9022_ (.CLK(clk),
    .D(_0324_),
    .RESET_B(net196),
    .Q(\mem[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9023_ (.CLK(clk),
    .D(_0325_),
    .RESET_B(net176),
    .Q(\mem[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9024_ (.CLK(clk),
    .D(_0326_),
    .RESET_B(net182),
    .Q(\mem[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9025_ (.CLK(clk),
    .D(_0327_),
    .RESET_B(net188),
    .Q(\mem[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9026_ (.CLK(clk),
    .D(_0328_),
    .RESET_B(net188),
    .Q(\mem[10][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9027_ (.CLK(clk),
    .D(_0329_),
    .RESET_B(net190),
    .Q(\mem[10][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9028_ (.CLK(clk),
    .D(_0330_),
    .RESET_B(net190),
    .Q(\mem[10][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9029_ (.CLK(clk),
    .D(_0331_),
    .RESET_B(net214),
    .Q(\mem[10][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9030_ (.CLK(clk),
    .D(_0332_),
    .RESET_B(net216),
    .Q(\mem[10][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9031_ (.CLK(clk),
    .D(_0333_),
    .RESET_B(net214),
    .Q(\mem[10][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9032_ (.CLK(clk),
    .D(_0334_),
    .RESET_B(net216),
    .Q(\mem[10][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9033_ (.CLK(clk),
    .D(_0335_),
    .RESET_B(net239),
    .Q(\mem[10][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9034_ (.CLK(clk),
    .D(_0336_),
    .RESET_B(net224),
    .Q(\mem[10][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9035_ (.CLK(clk),
    .D(_0337_),
    .RESET_B(net220),
    .Q(\mem[10][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9036_ (.CLK(clk),
    .D(_0338_),
    .RESET_B(net211),
    .Q(\mem[10][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9037_ (.CLK(clk),
    .D(_0339_),
    .RESET_B(net219),
    .Q(\mem[10][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9038_ (.CLK(clk),
    .D(_0340_),
    .RESET_B(net167),
    .Q(\mem[10][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9039_ (.CLK(clk),
    .D(_0341_),
    .RESET_B(net167),
    .Q(\mem[10][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9040_ (.CLK(clk),
    .D(_0342_),
    .RESET_B(net159),
    .Q(\mem[10][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9041_ (.CLK(clk),
    .D(_0343_),
    .RESET_B(net168),
    .Q(\mem[10][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9042_ (.CLK(clk),
    .D(_0344_),
    .RESET_B(net165),
    .Q(\mem[10][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9043_ (.CLK(clk),
    .D(_0345_),
    .RESET_B(net160),
    .Q(\mem[10][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9044_ (.CLK(clk),
    .D(_0346_),
    .RESET_B(net157),
    .Q(\mem[10][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9045_ (.CLK(clk),
    .D(_0347_),
    .RESET_B(net160),
    .Q(\mem[10][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9046_ (.CLK(clk),
    .D(_0348_),
    .RESET_B(net157),
    .Q(\mem[10][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9047_ (.CLK(clk),
    .D(_0349_),
    .RESET_B(net131),
    .Q(\mem[10][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9048_ (.CLK(clk),
    .D(_0350_),
    .RESET_B(net130),
    .Q(\mem[10][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9049_ (.CLK(clk),
    .D(_0351_),
    .RESET_B(net130),
    .Q(\mem[10][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9050_ (.CLK(clk),
    .D(_0352_),
    .RESET_B(net187),
    .Q(\mem[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9051_ (.CLK(clk),
    .D(_0353_),
    .RESET_B(net126),
    .Q(\mem[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9052_ (.CLK(clk),
    .D(_0354_),
    .RESET_B(net126),
    .Q(\mem[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9053_ (.CLK(clk),
    .D(_0355_),
    .RESET_B(net198),
    .Q(\mem[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9054_ (.CLK(clk),
    .D(_0356_),
    .RESET_B(net194),
    .Q(\mem[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9055_ (.CLK(clk),
    .D(_0357_),
    .RESET_B(net175),
    .Q(\mem[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9056_ (.CLK(clk),
    .D(_0358_),
    .RESET_B(net179),
    .Q(\mem[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9057_ (.CLK(clk),
    .D(_0359_),
    .RESET_B(net198),
    .Q(\mem[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9058_ (.CLK(clk),
    .D(_0360_),
    .RESET_B(net206),
    .Q(\mem[11][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9059_ (.CLK(clk),
    .D(_0361_),
    .RESET_B(net208),
    .Q(\mem[11][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9060_ (.CLK(clk),
    .D(_0362_),
    .RESET_B(net209),
    .Q(\mem[11][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9061_ (.CLK(clk),
    .D(_0363_),
    .RESET_B(net233),
    .Q(\mem[11][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9062_ (.CLK(clk),
    .D(_0364_),
    .RESET_B(net227),
    .Q(\mem[11][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9063_ (.CLK(clk),
    .D(_0365_),
    .RESET_B(net235),
    .Q(\mem[11][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9064_ (.CLK(clk),
    .D(_0366_),
    .RESET_B(net235),
    .Q(\mem[11][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9065_ (.CLK(clk),
    .D(_0367_),
    .RESET_B(net241),
    .Q(\mem[11][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9066_ (.CLK(clk),
    .D(_0368_),
    .RESET_B(net243),
    .Q(\mem[11][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9067_ (.CLK(clk),
    .D(_0369_),
    .RESET_B(net226),
    .Q(\mem[11][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9068_ (.CLK(clk),
    .D(_0370_),
    .RESET_B(net222),
    .Q(\mem[11][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9069_ (.CLK(clk),
    .D(_0371_),
    .RESET_B(net171),
    .Q(\mem[11][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9070_ (.CLK(clk),
    .D(_0372_),
    .RESET_B(net150),
    .Q(\mem[11][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9071_ (.CLK(clk),
    .D(_0373_),
    .RESET_B(net150),
    .Q(\mem[11][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9072_ (.CLK(clk),
    .D(_0374_),
    .RESET_B(net140),
    .Q(\mem[11][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9073_ (.CLK(clk),
    .D(_0375_),
    .RESET_B(net148),
    .Q(\mem[11][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9074_ (.CLK(clk),
    .D(_0376_),
    .RESET_B(net148),
    .Q(\mem[11][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9075_ (.CLK(clk),
    .D(_0377_),
    .RESET_B(net140),
    .Q(\mem[11][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9076_ (.CLK(clk),
    .D(_0378_),
    .RESET_B(net137),
    .Q(\mem[11][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9077_ (.CLK(clk),
    .D(_0379_),
    .RESET_B(net137),
    .Q(\mem[11][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9078_ (.CLK(clk),
    .D(_0380_),
    .RESET_B(net115),
    .Q(\mem[11][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9079_ (.CLK(clk),
    .D(_0381_),
    .RESET_B(net114),
    .Q(\mem[11][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9080_ (.CLK(clk),
    .D(_0382_),
    .RESET_B(net121),
    .Q(\mem[11][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9081_ (.CLK(clk),
    .D(_0383_),
    .RESET_B(net117),
    .Q(\mem[11][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9082_ (.CLK(clk),
    .D(_0384_),
    .RESET_B(net186),
    .Q(\mem[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9083_ (.CLK(clk),
    .D(_0385_),
    .RESET_B(net123),
    .Q(\mem[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9084_ (.CLK(clk),
    .D(_0386_),
    .RESET_B(net123),
    .Q(\mem[12][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9085_ (.CLK(clk),
    .D(_0387_),
    .RESET_B(net196),
    .Q(\mem[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9086_ (.CLK(clk),
    .D(_0388_),
    .RESET_B(net196),
    .Q(\mem[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9087_ (.CLK(clk),
    .D(_0389_),
    .RESET_B(net177),
    .Q(\mem[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9088_ (.CLK(clk),
    .D(_0390_),
    .RESET_B(net182),
    .Q(\mem[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9089_ (.CLK(clk),
    .D(_0391_),
    .RESET_B(net201),
    .Q(\mem[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9090_ (.CLK(clk),
    .D(_0392_),
    .RESET_B(net201),
    .Q(\mem[12][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9091_ (.CLK(clk),
    .D(_0393_),
    .RESET_B(net203),
    .Q(\mem[12][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9092_ (.CLK(clk),
    .D(_0394_),
    .RESET_B(net203),
    .Q(\mem[12][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9093_ (.CLK(clk),
    .D(_0395_),
    .RESET_B(net230),
    .Q(\mem[12][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9094_ (.CLK(clk),
    .D(_0396_),
    .RESET_B(net216),
    .Q(\mem[12][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9095_ (.CLK(clk),
    .D(_0397_),
    .RESET_B(net229),
    .Q(\mem[12][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9096_ (.CLK(clk),
    .D(_0398_),
    .RESET_B(net232),
    .Q(\mem[12][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9097_ (.CLK(clk),
    .D(_0399_),
    .RESET_B(net238),
    .Q(\mem[12][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9098_ (.CLK(clk),
    .D(_0400_),
    .RESET_B(net238),
    .Q(\mem[12][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9099_ (.CLK(clk),
    .D(_0401_),
    .RESET_B(net216),
    .Q(\mem[12][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9100_ (.CLK(clk),
    .D(_0402_),
    .RESET_B(net161),
    .Q(\mem[12][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9101_ (.CLK(clk),
    .D(_0403_),
    .RESET_B(net169),
    .Q(\mem[12][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9102_ (.CLK(clk),
    .D(_0404_),
    .RESET_B(net165),
    .Q(\mem[12][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9103_ (.CLK(clk),
    .D(_0405_),
    .RESET_B(net153),
    .Q(\mem[12][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9104_ (.CLK(clk),
    .D(_0406_),
    .RESET_B(net146),
    .Q(\mem[12][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9105_ (.CLK(clk),
    .D(_0407_),
    .RESET_B(net153),
    .Q(\mem[12][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9106_ (.CLK(clk),
    .D(_0408_),
    .RESET_B(net153),
    .Q(\mem[12][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9107_ (.CLK(clk),
    .D(_0409_),
    .RESET_B(net146),
    .Q(\mem[12][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9108_ (.CLK(clk),
    .D(_0410_),
    .RESET_B(net144),
    .Q(\mem[12][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9109_ (.CLK(clk),
    .D(_0411_),
    .RESET_B(net144),
    .Q(\mem[12][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9110_ (.CLK(clk),
    .D(_0412_),
    .RESET_B(net119),
    .Q(\mem[12][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9111_ (.CLK(clk),
    .D(_0413_),
    .RESET_B(net119),
    .Q(\mem[12][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9112_ (.CLK(clk),
    .D(_0414_),
    .RESET_B(net116),
    .Q(\mem[12][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9113_ (.CLK(clk),
    .D(_0415_),
    .RESET_B(net116),
    .Q(\mem[12][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9114_ (.CLK(clk),
    .D(_0416_),
    .RESET_B(net186),
    .Q(\mem[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9115_ (.CLK(clk),
    .D(_0417_),
    .RESET_B(net128),
    .Q(\mem[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9116_ (.CLK(clk),
    .D(_0418_),
    .RESET_B(net127),
    .Q(\mem[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9117_ (.CLK(clk),
    .D(_0419_),
    .RESET_B(net182),
    .Q(\mem[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9118_ (.CLK(clk),
    .D(_0420_),
    .RESET_B(net182),
    .Q(\mem[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9119_ (.CLK(clk),
    .D(_0421_),
    .RESET_B(net185),
    .Q(\mem[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9120_ (.CLK(clk),
    .D(_0422_),
    .RESET_B(net177),
    .Q(\mem[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9121_ (.CLK(clk),
    .D(_0423_),
    .RESET_B(net189),
    .Q(\mem[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9122_ (.CLK(clk),
    .D(_0424_),
    .RESET_B(net189),
    .Q(\mem[13][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9123_ (.CLK(clk),
    .D(_0425_),
    .RESET_B(net191),
    .Q(\mem[13][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9124_ (.CLK(clk),
    .D(_0426_),
    .RESET_B(net191),
    .Q(\mem[13][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9125_ (.CLK(clk),
    .D(_0427_),
    .RESET_B(net214),
    .Q(\mem[13][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9126_ (.CLK(clk),
    .D(_0428_),
    .RESET_B(net216),
    .Q(\mem[13][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9127_ (.CLK(clk),
    .D(_0429_),
    .RESET_B(net215),
    .Q(\mem[13][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9128_ (.CLK(clk),
    .D(_0430_),
    .RESET_B(net217),
    .Q(\mem[13][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9129_ (.CLK(clk),
    .D(_0431_),
    .RESET_B(net217),
    .Q(\mem[13][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9130_ (.CLK(clk),
    .D(_0432_),
    .RESET_B(net217),
    .Q(\mem[13][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9131_ (.CLK(clk),
    .D(_0433_),
    .RESET_B(net212),
    .Q(\mem[13][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9132_ (.CLK(clk),
    .D(_0434_),
    .RESET_B(net212),
    .Q(\mem[13][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9133_ (.CLK(clk),
    .D(_0435_),
    .RESET_B(net219),
    .Q(\mem[13][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9134_ (.CLK(clk),
    .D(_0436_),
    .RESET_B(net169),
    .Q(\mem[13][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9135_ (.CLK(clk),
    .D(_0437_),
    .RESET_B(net165),
    .Q(\mem[13][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9136_ (.CLK(clk),
    .D(_0438_),
    .RESET_B(net160),
    .Q(\mem[13][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9137_ (.CLK(clk),
    .D(_0439_),
    .RESET_B(net165),
    .Q(\mem[13][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9138_ (.CLK(clk),
    .D(_0440_),
    .RESET_B(net165),
    .Q(\mem[13][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9139_ (.CLK(clk),
    .D(_0441_),
    .RESET_B(net160),
    .Q(\mem[13][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9140_ (.CLK(clk),
    .D(_0442_),
    .RESET_B(net163),
    .Q(\mem[13][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9141_ (.CLK(clk),
    .D(_0443_),
    .RESET_B(net162),
    .Q(\mem[13][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9142_ (.CLK(clk),
    .D(_0444_),
    .RESET_B(net157),
    .Q(\mem[13][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9143_ (.CLK(clk),
    .D(_0445_),
    .RESET_B(net131),
    .Q(\mem[13][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9144_ (.CLK(clk),
    .D(_0446_),
    .RESET_B(net132),
    .Q(\mem[13][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9145_ (.CLK(clk),
    .D(_0447_),
    .RESET_B(net130),
    .Q(\mem[13][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9146_ (.CLK(clk),
    .D(_0448_),
    .RESET_B(net134),
    .Q(\mem[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9147_ (.CLK(clk),
    .D(_0449_),
    .RESET_B(net126),
    .Q(\mem[14][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9148_ (.CLK(clk),
    .D(_0450_),
    .RESET_B(net125),
    .Q(\mem[14][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9149_ (.CLK(clk),
    .D(_0451_),
    .RESET_B(net198),
    .Q(\mem[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9150_ (.CLK(clk),
    .D(_0452_),
    .RESET_B(net194),
    .Q(\mem[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9151_ (.CLK(clk),
    .D(_0453_),
    .RESET_B(net175),
    .Q(\mem[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9152_ (.CLK(clk),
    .D(_0454_),
    .RESET_B(net180),
    .Q(\mem[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9153_ (.CLK(clk),
    .D(_0455_),
    .RESET_B(net199),
    .Q(\mem[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9154_ (.CLK(clk),
    .D(_0456_),
    .RESET_B(net206),
    .Q(\mem[14][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9155_ (.CLK(clk),
    .D(_0457_),
    .RESET_B(net208),
    .Q(\mem[14][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9156_ (.CLK(clk),
    .D(_0458_),
    .RESET_B(net208),
    .Q(\mem[14][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9157_ (.CLK(clk),
    .D(_0459_),
    .RESET_B(net237),
    .Q(\mem[14][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9158_ (.CLK(clk),
    .D(_0460_),
    .RESET_B(net227),
    .Q(\mem[14][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9159_ (.CLK(clk),
    .D(_0461_),
    .RESET_B(net235),
    .Q(\mem[14][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9160_ (.CLK(clk),
    .D(_0462_),
    .RESET_B(net235),
    .Q(\mem[14][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9161_ (.CLK(clk),
    .D(_0463_),
    .RESET_B(net241),
    .Q(\mem[14][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9162_ (.CLK(clk),
    .D(_0464_),
    .RESET_B(net243),
    .Q(\mem[14][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9163_ (.CLK(clk),
    .D(_0465_),
    .RESET_B(net226),
    .Q(\mem[14][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9164_ (.CLK(clk),
    .D(_0466_),
    .RESET_B(net222),
    .Q(\mem[14][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9165_ (.CLK(clk),
    .D(_0467_),
    .RESET_B(net171),
    .Q(\mem[14][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9166_ (.CLK(clk),
    .D(_0468_),
    .RESET_B(net150),
    .Q(\mem[14][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9167_ (.CLK(clk),
    .D(_0469_),
    .RESET_B(net151),
    .Q(\mem[14][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9168_ (.CLK(clk),
    .D(_0470_),
    .RESET_B(net140),
    .Q(\mem[14][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9169_ (.CLK(clk),
    .D(_0471_),
    .RESET_B(net148),
    .Q(\mem[14][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9170_ (.CLK(clk),
    .D(_0472_),
    .RESET_B(net149),
    .Q(\mem[14][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9171_ (.CLK(clk),
    .D(_0473_),
    .RESET_B(net140),
    .Q(\mem[14][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9172_ (.CLK(clk),
    .D(_0474_),
    .RESET_B(net137),
    .Q(\mem[14][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9173_ (.CLK(clk),
    .D(_0475_),
    .RESET_B(net139),
    .Q(\mem[14][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9174_ (.CLK(clk),
    .D(_0476_),
    .RESET_B(net115),
    .Q(\mem[14][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9175_ (.CLK(clk),
    .D(_0477_),
    .RESET_B(net114),
    .Q(\mem[14][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9176_ (.CLK(clk),
    .D(_0478_),
    .RESET_B(net121),
    .Q(\mem[14][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9177_ (.CLK(clk),
    .D(_0479_),
    .RESET_B(net121),
    .Q(\mem[14][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9178_ (.CLK(clk),
    .D(_0480_),
    .RESET_B(net186),
    .Q(\mem[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9179_ (.CLK(clk),
    .D(_0481_),
    .RESET_B(net176),
    .Q(\mem[15][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9180_ (.CLK(clk),
    .D(_0482_),
    .RESET_B(net176),
    .Q(\mem[15][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9181_ (.CLK(clk),
    .D(_0483_),
    .RESET_B(net182),
    .Q(\mem[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9182_ (.CLK(clk),
    .D(_0484_),
    .RESET_B(net182),
    .Q(\mem[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9183_ (.CLK(clk),
    .D(_0485_),
    .RESET_B(net177),
    .Q(\mem[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9184_ (.CLK(clk),
    .D(_0486_),
    .RESET_B(net182),
    .Q(\mem[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9185_ (.CLK(clk),
    .D(_0487_),
    .RESET_B(net189),
    .Q(\mem[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9186_ (.CLK(clk),
    .D(_0488_),
    .RESET_B(net189),
    .Q(\mem[15][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9187_ (.CLK(clk),
    .D(_0489_),
    .RESET_B(net191),
    .Q(\mem[15][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9188_ (.CLK(clk),
    .D(_0490_),
    .RESET_B(net215),
    .Q(\mem[15][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9189_ (.CLK(clk),
    .D(_0491_),
    .RESET_B(net215),
    .Q(\mem[15][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9190_ (.CLK(clk),
    .D(_0492_),
    .RESET_B(net217),
    .Q(\mem[15][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9191_ (.CLK(clk),
    .D(_0493_),
    .RESET_B(net215),
    .Q(\mem[15][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9192_ (.CLK(clk),
    .D(_0494_),
    .RESET_B(net217),
    .Q(\mem[15][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9193_ (.CLK(clk),
    .D(_0495_),
    .RESET_B(net225),
    .Q(\mem[15][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9194_ (.CLK(clk),
    .D(_0496_),
    .RESET_B(net225),
    .Q(\mem[15][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9195_ (.CLK(clk),
    .D(_0497_),
    .RESET_B(net220),
    .Q(\mem[15][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9196_ (.CLK(clk),
    .D(_0498_),
    .RESET_B(net212),
    .Q(\mem[15][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9197_ (.CLK(clk),
    .D(_0499_),
    .RESET_B(net219),
    .Q(\mem[15][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9198_ (.CLK(clk),
    .D(_0500_),
    .RESET_B(net167),
    .Q(\mem[15][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9199_ (.CLK(clk),
    .D(_0501_),
    .RESET_B(net172),
    .Q(\mem[15][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9200_ (.CLK(clk),
    .D(_0502_),
    .RESET_B(net160),
    .Q(\mem[15][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9201_ (.CLK(clk),
    .D(_0503_),
    .RESET_B(net167),
    .Q(\mem[15][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9202_ (.CLK(clk),
    .D(_0504_),
    .RESET_B(net160),
    .Q(\mem[15][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9203_ (.CLK(clk),
    .D(_0505_),
    .RESET_B(net160),
    .Q(\mem[15][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9204_ (.CLK(clk),
    .D(_0506_),
    .RESET_B(net157),
    .Q(\mem[15][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9205_ (.CLK(clk),
    .D(_0507_),
    .RESET_B(net158),
    .Q(\mem[15][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9206_ (.CLK(clk),
    .D(_0508_),
    .RESET_B(net158),
    .Q(\mem[15][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9207_ (.CLK(clk),
    .D(_0509_),
    .RESET_B(net132),
    .Q(\mem[15][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9208_ (.CLK(clk),
    .D(_0510_),
    .RESET_B(net130),
    .Q(\mem[15][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9209_ (.CLK(clk),
    .D(_0511_),
    .RESET_B(net133),
    .Q(\mem[15][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9210_ (.CLK(clk),
    .D(_0512_),
    .RESET_B(net184),
    .Q(\mem[16][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9211_ (.CLK(clk),
    .D(_0513_),
    .RESET_B(net174),
    .Q(\mem[16][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9212_ (.CLK(clk),
    .D(_0514_),
    .RESET_B(net174),
    .Q(\mem[16][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9213_ (.CLK(clk),
    .D(_0515_),
    .RESET_B(net195),
    .Q(\mem[16][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9214_ (.CLK(clk),
    .D(_0516_),
    .RESET_B(net180),
    .Q(\mem[16][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9215_ (.CLK(clk),
    .D(_0517_),
    .RESET_B(net174),
    .Q(\mem[16][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9216_ (.CLK(clk),
    .D(_0518_),
    .RESET_B(net179),
    .Q(\mem[16][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9217_ (.CLK(clk),
    .D(_0519_),
    .RESET_B(net205),
    .Q(\mem[16][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9218_ (.CLK(clk),
    .D(_0520_),
    .RESET_B(net205),
    .Q(\mem[16][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9219_ (.CLK(clk),
    .D(_0521_),
    .RESET_B(net207),
    .Q(\mem[16][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9220_ (.CLK(clk),
    .D(_0522_),
    .RESET_B(net207),
    .Q(\mem[16][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9221_ (.CLK(clk),
    .D(_0523_),
    .RESET_B(net234),
    .Q(\mem[16][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9222_ (.CLK(clk),
    .D(_0524_),
    .RESET_B(net226),
    .Q(\mem[16][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9223_ (.CLK(clk),
    .D(_0525_),
    .RESET_B(net234),
    .Q(\mem[16][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9224_ (.CLK(clk),
    .D(_0526_),
    .RESET_B(net236),
    .Q(\mem[16][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9225_ (.CLK(clk),
    .D(_0527_),
    .RESET_B(net240),
    .Q(\mem[16][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9226_ (.CLK(clk),
    .D(_0528_),
    .RESET_B(net242),
    .Q(\mem[16][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9227_ (.CLK(clk),
    .D(_0529_),
    .RESET_B(net222),
    .Q(\mem[16][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9228_ (.CLK(clk),
    .D(_0530_),
    .RESET_B(net219),
    .Q(\mem[16][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9229_ (.CLK(clk),
    .D(_0531_),
    .RESET_B(net222),
    .Q(\mem[16][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9230_ (.CLK(clk),
    .D(_0532_),
    .RESET_B(net155),
    .Q(\mem[16][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9231_ (.CLK(clk),
    .D(_0533_),
    .RESET_B(net152),
    .Q(\mem[16][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9232_ (.CLK(clk),
    .D(_0534_),
    .RESET_B(net141),
    .Q(\mem[16][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9233_ (.CLK(clk),
    .D(_0535_),
    .RESET_B(net154),
    .Q(\mem[16][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9234_ (.CLK(clk),
    .D(_0536_),
    .RESET_B(net149),
    .Q(\mem[16][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9235_ (.CLK(clk),
    .D(_0537_),
    .RESET_B(net145),
    .Q(\mem[16][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9236_ (.CLK(clk),
    .D(_0538_),
    .RESET_B(net143),
    .Q(\mem[16][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9237_ (.CLK(clk),
    .D(_0539_),
    .RESET_B(net138),
    .Q(\mem[16][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9238_ (.CLK(clk),
    .D(_0540_),
    .RESET_B(net118),
    .Q(\mem[16][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9239_ (.CLK(clk),
    .D(_0541_),
    .RESET_B(net118),
    .Q(\mem[16][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9240_ (.CLK(clk),
    .D(_0542_),
    .RESET_B(net136),
    .Q(\mem[16][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9241_ (.CLK(clk),
    .D(_0543_),
    .RESET_B(net136),
    .Q(\mem[16][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9242_ (.CLK(clk),
    .D(_0544_),
    .RESET_B(net186),
    .Q(\mem[17][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9243_ (.CLK(clk),
    .D(_0545_),
    .RESET_B(net125),
    .Q(\mem[17][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9244_ (.CLK(clk),
    .D(_0546_),
    .RESET_B(net125),
    .Q(\mem[17][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9245_ (.CLK(clk),
    .D(_0547_),
    .RESET_B(net199),
    .Q(\mem[17][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9246_ (.CLK(clk),
    .D(_0548_),
    .RESET_B(net195),
    .Q(\mem[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9247_ (.CLK(clk),
    .D(_0549_),
    .RESET_B(net175),
    .Q(\mem[17][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9248_ (.CLK(clk),
    .D(_0550_),
    .RESET_B(net179),
    .Q(\mem[17][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9249_ (.CLK(clk),
    .D(_0551_),
    .RESET_B(net198),
    .Q(\mem[17][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9250_ (.CLK(clk),
    .D(_0552_),
    .RESET_B(net205),
    .Q(\mem[17][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9251_ (.CLK(clk),
    .D(_0553_),
    .RESET_B(net207),
    .Q(\mem[17][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9252_ (.CLK(clk),
    .D(_0554_),
    .RESET_B(net207),
    .Q(\mem[17][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9253_ (.CLK(clk),
    .D(_0555_),
    .RESET_B(net234),
    .Q(\mem[17][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9254_ (.CLK(clk),
    .D(_0556_),
    .RESET_B(net240),
    .Q(\mem[17][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9255_ (.CLK(clk),
    .D(_0557_),
    .RESET_B(net236),
    .Q(\mem[17][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9256_ (.CLK(clk),
    .D(_0558_),
    .RESET_B(net236),
    .Q(\mem[17][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9257_ (.CLK(clk),
    .D(_0559_),
    .RESET_B(net244),
    .Q(\mem[17][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9258_ (.CLK(clk),
    .D(_0560_),
    .RESET_B(net242),
    .Q(\mem[17][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9259_ (.CLK(clk),
    .D(_0561_),
    .RESET_B(net223),
    .Q(\mem[17][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9260_ (.CLK(clk),
    .D(_0562_),
    .RESET_B(net213),
    .Q(\mem[17][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9261_ (.CLK(clk),
    .D(_0563_),
    .RESET_B(net171),
    .Q(\mem[17][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9262_ (.CLK(clk),
    .D(_0564_),
    .RESET_B(net166),
    .Q(\mem[17][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9263_ (.CLK(clk),
    .D(_0565_),
    .RESET_B(net154),
    .Q(\mem[17][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9264_ (.CLK(clk),
    .D(_0566_),
    .RESET_B(net141),
    .Q(\mem[17][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9265_ (.CLK(clk),
    .D(_0567_),
    .RESET_B(net155),
    .Q(\mem[17][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9266_ (.CLK(clk),
    .D(_0568_),
    .RESET_B(net149),
    .Q(\mem[17][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9267_ (.CLK(clk),
    .D(_0569_),
    .RESET_B(net141),
    .Q(\mem[17][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9268_ (.CLK(clk),
    .D(_0570_),
    .RESET_B(net138),
    .Q(\mem[17][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9269_ (.CLK(clk),
    .D(_0571_),
    .RESET_B(net138),
    .Q(\mem[17][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9270_ (.CLK(clk),
    .D(_0572_),
    .RESET_B(net114),
    .Q(\mem[17][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9271_ (.CLK(clk),
    .D(_0573_),
    .RESET_B(net131),
    .Q(\mem[17][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9272_ (.CLK(clk),
    .D(_0574_),
    .RESET_B(net122),
    .Q(\mem[17][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9273_ (.CLK(clk),
    .D(_0575_),
    .RESET_B(net122),
    .Q(\mem[17][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9274_ (.CLK(clk),
    .D(_0576_),
    .RESET_B(net135),
    .Q(\mem[18][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9275_ (.CLK(clk),
    .D(_0577_),
    .RESET_B(net128),
    .Q(\mem[18][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9276_ (.CLK(clk),
    .D(_0578_),
    .RESET_B(net127),
    .Q(\mem[18][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9277_ (.CLK(clk),
    .D(_0579_),
    .RESET_B(net180),
    .Q(\mem[18][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9278_ (.CLK(clk),
    .D(_0580_),
    .RESET_B(net180),
    .Q(\mem[18][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9279_ (.CLK(clk),
    .D(_0581_),
    .RESET_B(net176),
    .Q(\mem[18][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9280_ (.CLK(clk),
    .D(_0582_),
    .RESET_B(net182),
    .Q(\mem[18][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9281_ (.CLK(clk),
    .D(_0583_),
    .RESET_B(net201),
    .Q(\mem[18][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9282_ (.CLK(clk),
    .D(_0584_),
    .RESET_B(net189),
    .Q(\mem[18][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9283_ (.CLK(clk),
    .D(_0585_),
    .RESET_B(net191),
    .Q(\mem[18][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9284_ (.CLK(clk),
    .D(_0586_),
    .RESET_B(net230),
    .Q(\mem[18][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9285_ (.CLK(clk),
    .D(_0587_),
    .RESET_B(net230),
    .Q(\mem[18][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9286_ (.CLK(clk),
    .D(_0588_),
    .RESET_B(net225),
    .Q(\mem[18][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9287_ (.CLK(clk),
    .D(_0589_),
    .RESET_B(net230),
    .Q(\mem[18][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9288_ (.CLK(clk),
    .D(_0590_),
    .RESET_B(net231),
    .Q(\mem[18][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9289_ (.CLK(clk),
    .D(_0591_),
    .RESET_B(net239),
    .Q(\mem[18][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9290_ (.CLK(clk),
    .D(_0592_),
    .RESET_B(net239),
    .Q(\mem[18][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9291_ (.CLK(clk),
    .D(_0593_),
    .RESET_B(net219),
    .Q(\mem[18][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9292_ (.CLK(clk),
    .D(_0594_),
    .RESET_B(net161),
    .Q(\mem[18][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9293_ (.CLK(clk),
    .D(_0595_),
    .RESET_B(net169),
    .Q(\mem[18][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9294_ (.CLK(clk),
    .D(_0596_),
    .RESET_B(net168),
    .Q(\mem[18][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9295_ (.CLK(clk),
    .D(_0597_),
    .RESET_B(net166),
    .Q(\mem[18][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9296_ (.CLK(clk),
    .D(_0598_),
    .RESET_B(net159),
    .Q(\mem[18][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9297_ (.CLK(clk),
    .D(_0599_),
    .RESET_B(net166),
    .Q(\mem[18][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9298_ (.CLK(clk),
    .D(_0600_),
    .RESET_B(net165),
    .Q(\mem[18][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9299_ (.CLK(clk),
    .D(_0601_),
    .RESET_B(net159),
    .Q(\mem[18][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9300_ (.CLK(clk),
    .D(_0602_),
    .RESET_B(net157),
    .Q(\mem[18][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9301_ (.CLK(clk),
    .D(_0603_),
    .RESET_B(net157),
    .Q(\mem[18][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9302_ (.CLK(clk),
    .D(_0604_),
    .RESET_B(net157),
    .Q(\mem[18][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9303_ (.CLK(clk),
    .D(_0605_),
    .RESET_B(net131),
    .Q(\mem[18][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9304_ (.CLK(clk),
    .D(_0606_),
    .RESET_B(net122),
    .Q(\mem[18][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9305_ (.CLK(clk),
    .D(_0607_),
    .RESET_B(net123),
    .Q(\mem[18][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9306_ (.CLK(clk),
    .D(_0608_),
    .RESET_B(net185),
    .Q(\mem[19][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9307_ (.CLK(clk),
    .D(_0609_),
    .RESET_B(net126),
    .Q(\mem[19][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9308_ (.CLK(clk),
    .D(_0610_),
    .RESET_B(net174),
    .Q(\mem[19][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9309_ (.CLK(clk),
    .D(_0611_),
    .RESET_B(net195),
    .Q(\mem[19][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9310_ (.CLK(clk),
    .D(_0612_),
    .RESET_B(net180),
    .Q(\mem[19][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9311_ (.CLK(clk),
    .D(_0613_),
    .RESET_B(net174),
    .Q(\mem[19][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9312_ (.CLK(clk),
    .D(_0614_),
    .RESET_B(net179),
    .Q(\mem[19][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9313_ (.CLK(clk),
    .D(_0615_),
    .RESET_B(net202),
    .Q(\mem[19][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9314_ (.CLK(clk),
    .D(_0616_),
    .RESET_B(net202),
    .Q(\mem[19][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9315_ (.CLK(clk),
    .D(_0617_),
    .RESET_B(net204),
    .Q(\mem[19][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9316_ (.CLK(clk),
    .D(_0618_),
    .RESET_B(net207),
    .Q(\mem[19][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9317_ (.CLK(clk),
    .D(_0619_),
    .RESET_B(net234),
    .Q(\mem[19][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9318_ (.CLK(clk),
    .D(_0620_),
    .RESET_B(net226),
    .Q(\mem[19][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9319_ (.CLK(clk),
    .D(_0621_),
    .RESET_B(net234),
    .Q(\mem[19][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9320_ (.CLK(clk),
    .D(_0622_),
    .RESET_B(net236),
    .Q(\mem[19][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9321_ (.CLK(clk),
    .D(_0623_),
    .RESET_B(net240),
    .Q(\mem[19][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9322_ (.CLK(clk),
    .D(_0624_),
    .RESET_B(net242),
    .Q(\mem[19][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9323_ (.CLK(clk),
    .D(_0625_),
    .RESET_B(net223),
    .Q(\mem[19][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9324_ (.CLK(clk),
    .D(_0626_),
    .RESET_B(net211),
    .Q(\mem[19][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9325_ (.CLK(clk),
    .D(_0627_),
    .RESET_B(net221),
    .Q(\mem[19][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9326_ (.CLK(clk),
    .D(_0628_),
    .RESET_B(net155),
    .Q(\mem[19][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9327_ (.CLK(clk),
    .D(_0629_),
    .RESET_B(net152),
    .Q(\mem[19][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9328_ (.CLK(clk),
    .D(_0630_),
    .RESET_B(net145),
    .Q(\mem[19][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9329_ (.CLK(clk),
    .D(_0631_),
    .RESET_B(net154),
    .Q(\mem[19][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9330_ (.CLK(clk),
    .D(_0632_),
    .RESET_B(net152),
    .Q(\mem[19][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9331_ (.CLK(clk),
    .D(_0633_),
    .RESET_B(net145),
    .Q(\mem[19][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9332_ (.CLK(clk),
    .D(_0634_),
    .RESET_B(net143),
    .Q(\mem[19][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9333_ (.CLK(clk),
    .D(_0635_),
    .RESET_B(net143),
    .Q(\mem[19][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9334_ (.CLK(clk),
    .D(_0636_),
    .RESET_B(net118),
    .Q(\mem[19][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9335_ (.CLK(clk),
    .D(_0637_),
    .RESET_B(net119),
    .Q(\mem[19][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9336_ (.CLK(clk),
    .D(_0638_),
    .RESET_B(net130),
    .Q(\mem[19][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9337_ (.CLK(clk),
    .D(_0639_),
    .RESET_B(net116),
    .Q(\mem[19][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9338_ (.CLK(clk),
    .D(_0640_),
    .RESET_B(net184),
    .Q(\mem[20][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9339_ (.CLK(clk),
    .D(_0641_),
    .RESET_B(net127),
    .Q(\mem[20][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9340_ (.CLK(clk),
    .D(_0642_),
    .RESET_B(net127),
    .Q(\mem[20][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9341_ (.CLK(clk),
    .D(_0643_),
    .RESET_B(net196),
    .Q(\mem[20][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9342_ (.CLK(clk),
    .D(_0644_),
    .RESET_B(net183),
    .Q(\mem[20][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9343_ (.CLK(clk),
    .D(_0645_),
    .RESET_B(net176),
    .Q(\mem[20][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9344_ (.CLK(clk),
    .D(_0646_),
    .RESET_B(net177),
    .Q(\mem[20][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9345_ (.CLK(clk),
    .D(_0647_),
    .RESET_B(net201),
    .Q(\mem[20][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9346_ (.CLK(clk),
    .D(_0648_),
    .RESET_B(net201),
    .Q(\mem[20][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9347_ (.CLK(clk),
    .D(_0649_),
    .RESET_B(net203),
    .Q(\mem[20][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9348_ (.CLK(clk),
    .D(_0650_),
    .RESET_B(net230),
    .Q(\mem[20][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9349_ (.CLK(clk),
    .D(_0651_),
    .RESET_B(net230),
    .Q(\mem[20][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9350_ (.CLK(clk),
    .D(_0652_),
    .RESET_B(net239),
    .Q(\mem[20][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9351_ (.CLK(clk),
    .D(_0653_),
    .RESET_B(net231),
    .Q(\mem[20][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9352_ (.CLK(clk),
    .D(_0654_),
    .RESET_B(net231),
    .Q(\mem[20][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9353_ (.CLK(clk),
    .D(_0655_),
    .RESET_B(net239),
    .Q(\mem[20][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9354_ (.CLK(clk),
    .D(_0656_),
    .RESET_B(net238),
    .Q(\mem[20][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9355_ (.CLK(clk),
    .D(_0657_),
    .RESET_B(net219),
    .Q(\mem[20][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9356_ (.CLK(clk),
    .D(_0658_),
    .RESET_B(net161),
    .Q(\mem[20][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9357_ (.CLK(clk),
    .D(_0659_),
    .RESET_B(net169),
    .Q(\mem[20][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9358_ (.CLK(clk),
    .D(_0660_),
    .RESET_B(net168),
    .Q(\mem[20][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9359_ (.CLK(clk),
    .D(_0661_),
    .RESET_B(net155),
    .Q(\mem[20][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9360_ (.CLK(clk),
    .D(_0662_),
    .RESET_B(net159),
    .Q(\mem[20][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9361_ (.CLK(clk),
    .D(_0663_),
    .RESET_B(net155),
    .Q(\mem[20][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9362_ (.CLK(clk),
    .D(_0664_),
    .RESET_B(net165),
    .Q(\mem[20][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9363_ (.CLK(clk),
    .D(_0665_),
    .RESET_B(net159),
    .Q(\mem[20][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9364_ (.CLK(clk),
    .D(_0666_),
    .RESET_B(net157),
    .Q(\mem[20][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9365_ (.CLK(clk),
    .D(_0667_),
    .RESET_B(net159),
    .Q(\mem[20][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9366_ (.CLK(clk),
    .D(_0668_),
    .RESET_B(net157),
    .Q(\mem[20][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9367_ (.CLK(clk),
    .D(_0669_),
    .RESET_B(net131),
    .Q(\mem[20][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9368_ (.CLK(clk),
    .D(_0670_),
    .RESET_B(net122),
    .Q(\mem[20][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9369_ (.CLK(clk),
    .D(_0671_),
    .RESET_B(net123),
    .Q(\mem[20][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9370_ (.CLK(clk),
    .D(_0672_),
    .RESET_B(net186),
    .Q(\mem[21][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9371_ (.CLK(clk),
    .D(_0673_),
    .RESET_B(net125),
    .Q(\mem[21][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9372_ (.CLK(clk),
    .D(_0674_),
    .RESET_B(net125),
    .Q(\mem[21][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9373_ (.CLK(clk),
    .D(_0675_),
    .RESET_B(net199),
    .Q(\mem[21][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9374_ (.CLK(clk),
    .D(_0676_),
    .RESET_B(net195),
    .Q(\mem[21][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9375_ (.CLK(clk),
    .D(_0677_),
    .RESET_B(net175),
    .Q(\mem[21][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9376_ (.CLK(clk),
    .D(_0678_),
    .RESET_B(net181),
    .Q(\mem[21][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9377_ (.CLK(clk),
    .D(_0679_),
    .RESET_B(net198),
    .Q(\mem[21][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9378_ (.CLK(clk),
    .D(_0680_),
    .RESET_B(net205),
    .Q(\mem[21][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9379_ (.CLK(clk),
    .D(_0681_),
    .RESET_B(net207),
    .Q(\mem[21][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9380_ (.CLK(clk),
    .D(_0682_),
    .RESET_B(net209),
    .Q(\mem[21][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9381_ (.CLK(clk),
    .D(_0683_),
    .RESET_B(net234),
    .Q(\mem[21][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9382_ (.CLK(clk),
    .D(_0684_),
    .RESET_B(net240),
    .Q(\mem[21][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9383_ (.CLK(clk),
    .D(_0685_),
    .RESET_B(net236),
    .Q(\mem[21][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9384_ (.CLK(clk),
    .D(_0686_),
    .RESET_B(net236),
    .Q(\mem[21][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9385_ (.CLK(clk),
    .D(_0687_),
    .RESET_B(net244),
    .Q(\mem[21][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9386_ (.CLK(clk),
    .D(_0688_),
    .RESET_B(net242),
    .Q(\mem[21][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9387_ (.CLK(clk),
    .D(_0689_),
    .RESET_B(net223),
    .Q(\mem[21][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9388_ (.CLK(clk),
    .D(_0690_),
    .RESET_B(net163),
    .Q(\mem[21][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9389_ (.CLK(clk),
    .D(_0691_),
    .RESET_B(net171),
    .Q(\mem[21][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9390_ (.CLK(clk),
    .D(_0692_),
    .RESET_B(net166),
    .Q(\mem[21][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9391_ (.CLK(clk),
    .D(_0693_),
    .RESET_B(net154),
    .Q(\mem[21][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9392_ (.CLK(clk),
    .D(_0694_),
    .RESET_B(net141),
    .Q(\mem[21][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9393_ (.CLK(clk),
    .D(_0695_),
    .RESET_B(net155),
    .Q(\mem[21][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9394_ (.CLK(clk),
    .D(_0696_),
    .RESET_B(net149),
    .Q(\mem[21][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9395_ (.CLK(clk),
    .D(_0697_),
    .RESET_B(net141),
    .Q(\mem[21][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9396_ (.CLK(clk),
    .D(_0698_),
    .RESET_B(net138),
    .Q(\mem[21][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9397_ (.CLK(clk),
    .D(_0699_),
    .RESET_B(net138),
    .Q(\mem[21][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9398_ (.CLK(clk),
    .D(_0700_),
    .RESET_B(net114),
    .Q(\mem[21][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9399_ (.CLK(clk),
    .D(_0701_),
    .RESET_B(net131),
    .Q(\mem[21][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9400_ (.CLK(clk),
    .D(_0702_),
    .RESET_B(net122),
    .Q(\mem[21][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9401_ (.CLK(clk),
    .D(_0703_),
    .RESET_B(net122),
    .Q(\mem[21][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9402_ (.CLK(clk),
    .D(_0704_),
    .RESET_B(net186),
    .Q(\mem[22][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9403_ (.CLK(clk),
    .D(_0705_),
    .RESET_B(net177),
    .Q(\mem[22][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9404_ (.CLK(clk),
    .D(_0706_),
    .RESET_B(net128),
    .Q(\mem[22][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9405_ (.CLK(clk),
    .D(_0707_),
    .RESET_B(net183),
    .Q(\mem[22][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9406_ (.CLK(clk),
    .D(_0708_),
    .RESET_B(net183),
    .Q(\mem[22][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9407_ (.CLK(clk),
    .D(_0709_),
    .RESET_B(net177),
    .Q(\mem[22][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9408_ (.CLK(clk),
    .D(_0710_),
    .RESET_B(net188),
    .Q(\mem[22][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9409_ (.CLK(clk),
    .D(_0711_),
    .RESET_B(net189),
    .Q(\mem[22][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9410_ (.CLK(clk),
    .D(_0712_),
    .RESET_B(net191),
    .Q(\mem[22][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9411_ (.CLK(clk),
    .D(_0713_),
    .RESET_B(net191),
    .Q(\mem[22][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9412_ (.CLK(clk),
    .D(_0714_),
    .RESET_B(net190),
    .Q(\mem[22][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9413_ (.CLK(clk),
    .D(_0715_),
    .RESET_B(net215),
    .Q(\mem[22][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9414_ (.CLK(clk),
    .D(_0716_),
    .RESET_B(net216),
    .Q(\mem[22][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9415_ (.CLK(clk),
    .D(_0717_),
    .RESET_B(net215),
    .Q(\mem[22][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9416_ (.CLK(clk),
    .D(_0718_),
    .RESET_B(net231),
    .Q(\mem[22][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9417_ (.CLK(clk),
    .D(_0719_),
    .RESET_B(net231),
    .Q(\mem[22][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9418_ (.CLK(clk),
    .D(_0720_),
    .RESET_B(net225),
    .Q(\mem[22][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9419_ (.CLK(clk),
    .D(_0721_),
    .RESET_B(net219),
    .Q(\mem[22][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9420_ (.CLK(clk),
    .D(_0722_),
    .RESET_B(net211),
    .Q(\mem[22][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9421_ (.CLK(clk),
    .D(_0723_),
    .RESET_B(net161),
    .Q(\mem[22][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9422_ (.CLK(clk),
    .D(_0724_),
    .RESET_B(net167),
    .Q(\mem[22][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9423_ (.CLK(clk),
    .D(_0725_),
    .RESET_B(net167),
    .Q(\mem[22][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9424_ (.CLK(clk),
    .D(_0726_),
    .RESET_B(net159),
    .Q(\mem[22][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9425_ (.CLK(clk),
    .D(_0727_),
    .RESET_B(net167),
    .Q(\mem[22][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9426_ (.CLK(clk),
    .D(_0728_),
    .RESET_B(net159),
    .Q(\mem[22][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9427_ (.CLK(clk),
    .D(_0729_),
    .RESET_B(net159),
    .Q(\mem[22][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9428_ (.CLK(clk),
    .D(_0730_),
    .RESET_B(net158),
    .Q(\mem[22][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9429_ (.CLK(clk),
    .D(_0731_),
    .RESET_B(net158),
    .Q(\mem[22][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9430_ (.CLK(clk),
    .D(_0732_),
    .RESET_B(net132),
    .Q(\mem[22][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9431_ (.CLK(clk),
    .D(_0733_),
    .RESET_B(net132),
    .Q(\mem[22][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9432_ (.CLK(clk),
    .D(_0734_),
    .RESET_B(net123),
    .Q(\mem[22][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9433_ (.CLK(clk),
    .D(_0735_),
    .RESET_B(net123),
    .Q(\mem[22][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9434_ (.CLK(clk),
    .D(_0736_),
    .RESET_B(net134),
    .Q(\mem[23][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9435_ (.CLK(clk),
    .D(_0737_),
    .RESET_B(net128),
    .Q(\mem[23][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9436_ (.CLK(clk),
    .D(_0738_),
    .RESET_B(net129),
    .Q(\mem[23][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9437_ (.CLK(clk),
    .D(_0739_),
    .RESET_B(net196),
    .Q(\mem[23][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9438_ (.CLK(clk),
    .D(_0740_),
    .RESET_B(net180),
    .Q(\mem[23][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9439_ (.CLK(clk),
    .D(_0741_),
    .RESET_B(net176),
    .Q(\mem[23][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9440_ (.CLK(clk),
    .D(_0742_),
    .RESET_B(net177),
    .Q(\mem[23][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9441_ (.CLK(clk),
    .D(_0743_),
    .RESET_B(net196),
    .Q(\mem[23][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9442_ (.CLK(clk),
    .D(_0744_),
    .RESET_B(net201),
    .Q(\mem[23][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9443_ (.CLK(clk),
    .D(_0745_),
    .RESET_B(net203),
    .Q(\mem[23][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9444_ (.CLK(clk),
    .D(_0746_),
    .RESET_B(net229),
    .Q(\mem[23][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9445_ (.CLK(clk),
    .D(_0747_),
    .RESET_B(net229),
    .Q(\mem[23][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9446_ (.CLK(clk),
    .D(_0748_),
    .RESET_B(net225),
    .Q(\mem[23][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9447_ (.CLK(clk),
    .D(_0749_),
    .RESET_B(net232),
    .Q(\mem[23][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9448_ (.CLK(clk),
    .D(_0750_),
    .RESET_B(net232),
    .Q(\mem[23][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9449_ (.CLK(clk),
    .D(_0751_),
    .RESET_B(net239),
    .Q(\mem[23][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9450_ (.CLK(clk),
    .D(_0752_),
    .RESET_B(net238),
    .Q(\mem[23][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9451_ (.CLK(clk),
    .D(_0753_),
    .RESET_B(net220),
    .Q(\mem[23][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9452_ (.CLK(clk),
    .D(_0754_),
    .RESET_B(net211),
    .Q(\mem[23][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9453_ (.CLK(clk),
    .D(_0755_),
    .RESET_B(net171),
    .Q(\mem[23][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9454_ (.CLK(clk),
    .D(_0756_),
    .RESET_B(net166),
    .Q(\mem[23][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9455_ (.CLK(clk),
    .D(_0757_),
    .RESET_B(net154),
    .Q(\mem[23][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9456_ (.CLK(clk),
    .D(_0758_),
    .RESET_B(net146),
    .Q(\mem[23][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9457_ (.CLK(clk),
    .D(_0759_),
    .RESET_B(net155),
    .Q(\mem[23][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9458_ (.CLK(clk),
    .D(_0760_),
    .RESET_B(net152),
    .Q(\mem[23][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9459_ (.CLK(clk),
    .D(_0761_),
    .RESET_B(net146),
    .Q(\mem[23][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9460_ (.CLK(clk),
    .D(_0762_),
    .RESET_B(net144),
    .Q(\mem[23][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9461_ (.CLK(clk),
    .D(_0763_),
    .RESET_B(net144),
    .Q(\mem[23][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9462_ (.CLK(clk),
    .D(_0764_),
    .RESET_B(net144),
    .Q(\mem[23][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9463_ (.CLK(clk),
    .D(_0765_),
    .RESET_B(net131),
    .Q(\mem[23][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9464_ (.CLK(clk),
    .D(_0766_),
    .RESET_B(net130),
    .Q(\mem[23][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9465_ (.CLK(clk),
    .D(_0767_),
    .RESET_B(net133),
    .Q(\mem[23][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9466_ (.CLK(clk),
    .D(_0768_),
    .RESET_B(net134),
    .Q(\mem[24][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9467_ (.CLK(clk),
    .D(_0769_),
    .RESET_B(net127),
    .Q(\mem[24][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9468_ (.CLK(clk),
    .D(_0770_),
    .RESET_B(net127),
    .Q(\mem[24][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9469_ (.CLK(clk),
    .D(_0771_),
    .RESET_B(net183),
    .Q(\mem[24][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9470_ (.CLK(clk),
    .D(_0772_),
    .RESET_B(net183),
    .Q(\mem[24][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9471_ (.CLK(clk),
    .D(_0773_),
    .RESET_B(net178),
    .Q(\mem[24][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9472_ (.CLK(clk),
    .D(_0774_),
    .RESET_B(net182),
    .Q(\mem[24][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9473_ (.CLK(clk),
    .D(_0775_),
    .RESET_B(net189),
    .Q(\mem[24][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9474_ (.CLK(clk),
    .D(_0776_),
    .RESET_B(net191),
    .Q(\mem[24][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9475_ (.CLK(clk),
    .D(_0777_),
    .RESET_B(net191),
    .Q(\mem[24][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9476_ (.CLK(clk),
    .D(_0778_),
    .RESET_B(net203),
    .Q(\mem[24][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9477_ (.CLK(clk),
    .D(_0779_),
    .RESET_B(net215),
    .Q(\mem[24][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9478_ (.CLK(clk),
    .D(_0780_),
    .RESET_B(net216),
    .Q(\mem[24][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9479_ (.CLK(clk),
    .D(_0781_),
    .RESET_B(net230),
    .Q(\mem[24][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9480_ (.CLK(clk),
    .D(_0782_),
    .RESET_B(net231),
    .Q(\mem[24][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9481_ (.CLK(clk),
    .D(_0783_),
    .RESET_B(net231),
    .Q(\mem[24][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9482_ (.CLK(clk),
    .D(_0784_),
    .RESET_B(net239),
    .Q(\mem[24][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9483_ (.CLK(clk),
    .D(_0785_),
    .RESET_B(net212),
    .Q(\mem[24][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9484_ (.CLK(clk),
    .D(_0786_),
    .RESET_B(net161),
    .Q(\mem[24][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9485_ (.CLK(clk),
    .D(_0787_),
    .RESET_B(net169),
    .Q(\mem[24][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9486_ (.CLK(clk),
    .D(_0788_),
    .RESET_B(net167),
    .Q(\mem[24][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9487_ (.CLK(clk),
    .D(_0789_),
    .RESET_B(net172),
    .Q(\mem[24][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9488_ (.CLK(clk),
    .D(_0790_),
    .RESET_B(net159),
    .Q(\mem[24][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9489_ (.CLK(clk),
    .D(_0791_),
    .RESET_B(net167),
    .Q(\mem[24][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9490_ (.CLK(clk),
    .D(_0792_),
    .RESET_B(net165),
    .Q(\mem[24][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9491_ (.CLK(clk),
    .D(_0793_),
    .RESET_B(net160),
    .Q(\mem[24][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9492_ (.CLK(clk),
    .D(_0794_),
    .RESET_B(net157),
    .Q(\mem[24][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9493_ (.CLK(clk),
    .D(_0795_),
    .RESET_B(net158),
    .Q(\mem[24][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9494_ (.CLK(clk),
    .D(_0796_),
    .RESET_B(net132),
    .Q(\mem[24][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9495_ (.CLK(clk),
    .D(_0797_),
    .RESET_B(net132),
    .Q(\mem[24][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9496_ (.CLK(clk),
    .D(_0798_),
    .RESET_B(net133),
    .Q(\mem[24][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9497_ (.CLK(clk),
    .D(_0799_),
    .RESET_B(net133),
    .Q(\mem[24][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9498_ (.CLK(clk),
    .D(_0800_),
    .RESET_B(net135),
    .Q(\mem[25][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9499_ (.CLK(clk),
    .D(_0801_),
    .RESET_B(net124),
    .Q(\mem[25][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9500_ (.CLK(clk),
    .D(_0802_),
    .RESET_B(net125),
    .Q(\mem[25][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9501_ (.CLK(clk),
    .D(_0803_),
    .RESET_B(net198),
    .Q(\mem[25][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9502_ (.CLK(clk),
    .D(_0804_),
    .RESET_B(net194),
    .Q(\mem[25][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9503_ (.CLK(clk),
    .D(_0805_),
    .RESET_B(net175),
    .Q(\mem[25][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9504_ (.CLK(clk),
    .D(_0806_),
    .RESET_B(net180),
    .Q(\mem[25][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9505_ (.CLK(clk),
    .D(_0807_),
    .RESET_B(net205),
    .Q(\mem[25][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9506_ (.CLK(clk),
    .D(_0808_),
    .RESET_B(net205),
    .Q(\mem[25][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9507_ (.CLK(clk),
    .D(_0809_),
    .RESET_B(net207),
    .Q(\mem[25][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9508_ (.CLK(clk),
    .D(_0810_),
    .RESET_B(net209),
    .Q(\mem[25][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9509_ (.CLK(clk),
    .D(_0811_),
    .RESET_B(net233),
    .Q(\mem[25][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9510_ (.CLK(clk),
    .D(_0812_),
    .RESET_B(net240),
    .Q(\mem[25][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9511_ (.CLK(clk),
    .D(_0813_),
    .RESET_B(net236),
    .Q(\mem[25][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9512_ (.CLK(clk),
    .D(_0814_),
    .RESET_B(net235),
    .Q(\mem[25][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9513_ (.CLK(clk),
    .D(_0815_),
    .RESET_B(net241),
    .Q(\mem[25][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9514_ (.CLK(clk),
    .D(_0816_),
    .RESET_B(net242),
    .Q(\mem[25][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9515_ (.CLK(clk),
    .D(_0817_),
    .RESET_B(net223),
    .Q(\mem[25][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9516_ (.CLK(clk),
    .D(_0818_),
    .RESET_B(net221),
    .Q(\mem[25][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9517_ (.CLK(clk),
    .D(_0819_),
    .RESET_B(net171),
    .Q(\mem[25][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9518_ (.CLK(clk),
    .D(_0820_),
    .RESET_B(net166),
    .Q(\mem[25][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9519_ (.CLK(clk),
    .D(_0821_),
    .RESET_B(net149),
    .Q(\mem[25][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9520_ (.CLK(clk),
    .D(_0822_),
    .RESET_B(net141),
    .Q(\mem[25][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9521_ (.CLK(clk),
    .D(_0823_),
    .RESET_B(net149),
    .Q(\mem[25][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9522_ (.CLK(clk),
    .D(_0824_),
    .RESET_B(net148),
    .Q(\mem[25][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9523_ (.CLK(clk),
    .D(_0825_),
    .RESET_B(net141),
    .Q(\mem[25][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9524_ (.CLK(clk),
    .D(_0826_),
    .RESET_B(net138),
    .Q(\mem[25][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9525_ (.CLK(clk),
    .D(_0827_),
    .RESET_B(net139),
    .Q(\mem[25][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9526_ (.CLK(clk),
    .D(_0828_),
    .RESET_B(net114),
    .Q(\mem[25][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9527_ (.CLK(clk),
    .D(_0829_),
    .RESET_B(net118),
    .Q(\mem[25][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9528_ (.CLK(clk),
    .D(_0830_),
    .RESET_B(net117),
    .Q(\mem[25][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9529_ (.CLK(clk),
    .D(_0831_),
    .RESET_B(net117),
    .Q(\mem[25][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9530_ (.CLK(clk),
    .D(_0832_),
    .RESET_B(net184),
    .Q(\mem[26][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9531_ (.CLK(clk),
    .D(_0833_),
    .RESET_B(net129),
    .Q(\mem[26][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9532_ (.CLK(clk),
    .D(_0834_),
    .RESET_B(net125),
    .Q(\mem[26][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9533_ (.CLK(clk),
    .D(_0835_),
    .RESET_B(net198),
    .Q(\mem[26][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9534_ (.CLK(clk),
    .D(_0836_),
    .RESET_B(net195),
    .Q(\mem[26][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9535_ (.CLK(clk),
    .D(_0837_),
    .RESET_B(net175),
    .Q(\mem[26][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9536_ (.CLK(clk),
    .D(_0838_),
    .RESET_B(net179),
    .Q(\mem[26][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9537_ (.CLK(clk),
    .D(_0839_),
    .RESET_B(net205),
    .Q(\mem[26][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9538_ (.CLK(clk),
    .D(_0840_),
    .RESET_B(net205),
    .Q(\mem[26][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9539_ (.CLK(clk),
    .D(_0841_),
    .RESET_B(net207),
    .Q(\mem[26][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9540_ (.CLK(clk),
    .D(_0842_),
    .RESET_B(net209),
    .Q(\mem[26][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9541_ (.CLK(clk),
    .D(_0843_),
    .RESET_B(net233),
    .Q(\mem[26][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9542_ (.CLK(clk),
    .D(_0844_),
    .RESET_B(net227),
    .Q(\mem[26][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9543_ (.CLK(clk),
    .D(_0845_),
    .RESET_B(net235),
    .Q(\mem[26][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9544_ (.CLK(clk),
    .D(_0846_),
    .RESET_B(net237),
    .Q(\mem[26][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9545_ (.CLK(clk),
    .D(_0847_),
    .RESET_B(net241),
    .Q(\mem[26][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9546_ (.CLK(clk),
    .D(_0848_),
    .RESET_B(net242),
    .Q(\mem[26][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9547_ (.CLK(clk),
    .D(_0849_),
    .RESET_B(net227),
    .Q(\mem[26][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9548_ (.CLK(clk),
    .D(_0850_),
    .RESET_B(net221),
    .Q(\mem[26][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9549_ (.CLK(clk),
    .D(_0851_),
    .RESET_B(net171),
    .Q(\mem[26][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9550_ (.CLK(clk),
    .D(_0852_),
    .RESET_B(net166),
    .Q(\mem[26][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9551_ (.CLK(clk),
    .D(_0853_),
    .RESET_B(net151),
    .Q(\mem[26][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9552_ (.CLK(clk),
    .D(_0854_),
    .RESET_B(net148),
    .Q(\mem[26][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9553_ (.CLK(clk),
    .D(_0855_),
    .RESET_B(net150),
    .Q(\mem[26][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9554_ (.CLK(clk),
    .D(_0856_),
    .RESET_B(net149),
    .Q(\mem[26][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9555_ (.CLK(clk),
    .D(_0857_),
    .RESET_B(net142),
    .Q(\mem[26][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9556_ (.CLK(clk),
    .D(_0858_),
    .RESET_B(net137),
    .Q(\mem[26][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9557_ (.CLK(clk),
    .D(_0859_),
    .RESET_B(net140),
    .Q(\mem[26][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9558_ (.CLK(clk),
    .D(_0860_),
    .RESET_B(net115),
    .Q(\mem[26][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9559_ (.CLK(clk),
    .D(_0861_),
    .RESET_B(net118),
    .Q(\mem[26][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9560_ (.CLK(clk),
    .D(_0862_),
    .RESET_B(net117),
    .Q(\mem[26][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9561_ (.CLK(clk),
    .D(_0863_),
    .RESET_B(net117),
    .Q(\mem[26][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9562_ (.CLK(clk),
    .D(_0864_),
    .RESET_B(net135),
    .Q(\mem[27][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9563_ (.CLK(clk),
    .D(_0865_),
    .RESET_B(net125),
    .Q(\mem[27][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9564_ (.CLK(clk),
    .D(_0866_),
    .RESET_B(net126),
    .Q(\mem[27][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9565_ (.CLK(clk),
    .D(_0867_),
    .RESET_B(net198),
    .Q(\mem[27][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9566_ (.CLK(clk),
    .D(_0868_),
    .RESET_B(net194),
    .Q(\mem[27][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9567_ (.CLK(clk),
    .D(_0869_),
    .RESET_B(net178),
    .Q(\mem[27][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9568_ (.CLK(clk),
    .D(_0870_),
    .RESET_B(net181),
    .Q(\mem[27][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9569_ (.CLK(clk),
    .D(_0871_),
    .RESET_B(net199),
    .Q(\mem[27][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9570_ (.CLK(clk),
    .D(_0872_),
    .RESET_B(net206),
    .Q(\mem[27][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9571_ (.CLK(clk),
    .D(_0873_),
    .RESET_B(net208),
    .Q(\mem[27][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9572_ (.CLK(clk),
    .D(_0874_),
    .RESET_B(net209),
    .Q(\mem[27][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9573_ (.CLK(clk),
    .D(_0875_),
    .RESET_B(net233),
    .Q(\mem[27][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9574_ (.CLK(clk),
    .D(_0876_),
    .RESET_B(net227),
    .Q(\mem[27][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9575_ (.CLK(clk),
    .D(_0877_),
    .RESET_B(net237),
    .Q(\mem[27][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9576_ (.CLK(clk),
    .D(_0878_),
    .RESET_B(net237),
    .Q(\mem[27][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9577_ (.CLK(clk),
    .D(_0879_),
    .RESET_B(net239),
    .Q(\mem[27][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9578_ (.CLK(clk),
    .D(_0880_),
    .RESET_B(net243),
    .Q(\mem[27][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9579_ (.CLK(clk),
    .D(_0881_),
    .RESET_B(net226),
    .Q(\mem[27][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9580_ (.CLK(clk),
    .D(_0882_),
    .RESET_B(net211),
    .Q(\mem[27][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9581_ (.CLK(clk),
    .D(_0883_),
    .RESET_B(net171),
    .Q(\mem[27][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9582_ (.CLK(clk),
    .D(_0884_),
    .RESET_B(net156),
    .Q(\mem[27][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9583_ (.CLK(clk),
    .D(_0885_),
    .RESET_B(net154),
    .Q(\mem[27][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9584_ (.CLK(clk),
    .D(_0886_),
    .RESET_B(net141),
    .Q(\mem[27][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9585_ (.CLK(clk),
    .D(_0887_),
    .RESET_B(net156),
    .Q(\mem[27][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9586_ (.CLK(clk),
    .D(_0888_),
    .RESET_B(net149),
    .Q(\mem[27][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9587_ (.CLK(clk),
    .D(_0889_),
    .RESET_B(net141),
    .Q(\mem[27][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9588_ (.CLK(clk),
    .D(_0890_),
    .RESET_B(net138),
    .Q(\mem[27][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9589_ (.CLK(clk),
    .D(_0891_),
    .RESET_B(net138),
    .Q(\mem[27][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9590_ (.CLK(clk),
    .D(_0892_),
    .RESET_B(net114),
    .Q(\mem[27][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9591_ (.CLK(clk),
    .D(_0893_),
    .RESET_B(net118),
    .Q(\mem[27][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9592_ (.CLK(clk),
    .D(_0894_),
    .RESET_B(net116),
    .Q(\mem[27][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9593_ (.CLK(clk),
    .D(_0895_),
    .RESET_B(net116),
    .Q(\mem[27][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9594_ (.CLK(clk),
    .D(_0896_),
    .RESET_B(net187),
    .Q(\mem[28][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9595_ (.CLK(clk),
    .D(_0897_),
    .RESET_B(net126),
    .Q(\mem[28][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9596_ (.CLK(clk),
    .D(_0898_),
    .RESET_B(net126),
    .Q(\mem[28][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9597_ (.CLK(clk),
    .D(_0899_),
    .RESET_B(net198),
    .Q(\mem[28][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9598_ (.CLK(clk),
    .D(_0900_),
    .RESET_B(net195),
    .Q(\mem[28][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9599_ (.CLK(clk),
    .D(_0901_),
    .RESET_B(net178),
    .Q(\mem[28][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9600_ (.CLK(clk),
    .D(_0902_),
    .RESET_B(net181),
    .Q(\mem[28][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9601_ (.CLK(clk),
    .D(_0903_),
    .RESET_B(net199),
    .Q(\mem[28][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9602_ (.CLK(clk),
    .D(_0904_),
    .RESET_B(net205),
    .Q(\mem[28][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9603_ (.CLK(clk),
    .D(_0905_),
    .RESET_B(net207),
    .Q(\mem[28][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9604_ (.CLK(clk),
    .D(_0906_),
    .RESET_B(net209),
    .Q(\mem[28][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9605_ (.CLK(clk),
    .D(_0907_),
    .RESET_B(net233),
    .Q(\mem[28][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9606_ (.CLK(clk),
    .D(_0908_),
    .RESET_B(net226),
    .Q(\mem[28][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9607_ (.CLK(clk),
    .D(_0909_),
    .RESET_B(net237),
    .Q(\mem[28][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9608_ (.CLK(clk),
    .D(_0910_),
    .RESET_B(net236),
    .Q(\mem[28][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9609_ (.CLK(clk),
    .D(_0911_),
    .RESET_B(net242),
    .Q(\mem[28][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9610_ (.CLK(clk),
    .D(_0912_),
    .RESET_B(net242),
    .Q(\mem[28][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9611_ (.CLK(clk),
    .D(_0913_),
    .RESET_B(net224),
    .Q(\mem[28][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9612_ (.CLK(clk),
    .D(_0914_),
    .RESET_B(net213),
    .Q(\mem[28][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9613_ (.CLK(clk),
    .D(_0915_),
    .RESET_B(net169),
    .Q(\mem[28][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9614_ (.CLK(clk),
    .D(_0916_),
    .RESET_B(net168),
    .Q(\mem[28][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9615_ (.CLK(clk),
    .D(_0917_),
    .RESET_B(net156),
    .Q(\mem[28][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9616_ (.CLK(clk),
    .D(_0918_),
    .RESET_B(net142),
    .Q(\mem[28][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9617_ (.CLK(clk),
    .D(_0919_),
    .RESET_B(net156),
    .Q(\mem[28][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9618_ (.CLK(clk),
    .D(_0920_),
    .RESET_B(net151),
    .Q(\mem[28][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9619_ (.CLK(clk),
    .D(_0921_),
    .RESET_B(net141),
    .Q(\mem[28][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9620_ (.CLK(clk),
    .D(_0922_),
    .RESET_B(net138),
    .Q(\mem[28][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9621_ (.CLK(clk),
    .D(_0923_),
    .RESET_B(net138),
    .Q(\mem[28][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9622_ (.CLK(clk),
    .D(_0924_),
    .RESET_B(net114),
    .Q(\mem[28][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9623_ (.CLK(clk),
    .D(_0925_),
    .RESET_B(net118),
    .Q(\mem[28][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9624_ (.CLK(clk),
    .D(_0926_),
    .RESET_B(net116),
    .Q(\mem[28][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9625_ (.CLK(clk),
    .D(_0927_),
    .RESET_B(net116),
    .Q(\mem[28][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9626_ (.CLK(clk),
    .D(_0928_),
    .RESET_B(net187),
    .Q(\mem[29][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9627_ (.CLK(clk),
    .D(_0929_),
    .RESET_B(net123),
    .Q(\mem[29][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9628_ (.CLK(clk),
    .D(_0930_),
    .RESET_B(net124),
    .Q(\mem[29][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9629_ (.CLK(clk),
    .D(_0931_),
    .RESET_B(net197),
    .Q(\mem[29][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9630_ (.CLK(clk),
    .D(_0932_),
    .RESET_B(net194),
    .Q(\mem[29][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9631_ (.CLK(clk),
    .D(_0933_),
    .RESET_B(net178),
    .Q(\mem[29][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9632_ (.CLK(clk),
    .D(_0934_),
    .RESET_B(net181),
    .Q(\mem[29][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9633_ (.CLK(clk),
    .D(_0935_),
    .RESET_B(net197),
    .Q(\mem[29][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9634_ (.CLK(clk),
    .D(_0936_),
    .RESET_B(net202),
    .Q(\mem[29][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9635_ (.CLK(clk),
    .D(_0937_),
    .RESET_B(net207),
    .Q(\mem[29][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9636_ (.CLK(clk),
    .D(_0938_),
    .RESET_B(net204),
    .Q(\mem[29][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9637_ (.CLK(clk),
    .D(_0939_),
    .RESET_B(net229),
    .Q(\mem[29][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9638_ (.CLK(clk),
    .D(_0940_),
    .RESET_B(net225),
    .Q(\mem[29][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9639_ (.CLK(clk),
    .D(_0941_),
    .RESET_B(net230),
    .Q(\mem[29][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9640_ (.CLK(clk),
    .D(_0942_),
    .RESET_B(net232),
    .Q(\mem[29][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9641_ (.CLK(clk),
    .D(_0943_),
    .RESET_B(net239),
    .Q(\mem[29][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9642_ (.CLK(clk),
    .D(_0944_),
    .RESET_B(net238),
    .Q(\mem[29][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9643_ (.CLK(clk),
    .D(_0945_),
    .RESET_B(net224),
    .Q(\mem[29][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9644_ (.CLK(clk),
    .D(_0946_),
    .RESET_B(net213),
    .Q(\mem[29][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9645_ (.CLK(clk),
    .D(_0947_),
    .RESET_B(net172),
    .Q(\mem[29][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9646_ (.CLK(clk),
    .D(_0948_),
    .RESET_B(net165),
    .Q(\mem[29][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9647_ (.CLK(clk),
    .D(_0949_),
    .RESET_B(net152),
    .Q(\mem[29][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9648_ (.CLK(clk),
    .D(_0950_),
    .RESET_B(net142),
    .Q(\mem[29][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9649_ (.CLK(clk),
    .D(_0951_),
    .RESET_B(net153),
    .Q(\mem[29][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9650_ (.CLK(clk),
    .D(_0952_),
    .RESET_B(net151),
    .Q(\mem[29][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9651_ (.CLK(clk),
    .D(_0953_),
    .RESET_B(net146),
    .Q(\mem[29][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9652_ (.CLK(clk),
    .D(_0954_),
    .RESET_B(net139),
    .Q(\mem[29][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9653_ (.CLK(clk),
    .D(_0955_),
    .RESET_B(net139),
    .Q(\mem[29][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9654_ (.CLK(clk),
    .D(_0956_),
    .RESET_B(net115),
    .Q(\mem[29][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9655_ (.CLK(clk),
    .D(_0957_),
    .RESET_B(net119),
    .Q(\mem[29][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9656_ (.CLK(clk),
    .D(_0958_),
    .RESET_B(net116),
    .Q(\mem[29][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9657_ (.CLK(clk),
    .D(_0959_),
    .RESET_B(net116),
    .Q(\mem[29][31] ));
 sky130_fd_sc_hd__dfrtp_1 _9658_ (.CLK(clk),
    .D(_0960_),
    .RESET_B(net187),
    .Q(\mem[30][0] ));
 sky130_fd_sc_hd__dfrtp_1 _9659_ (.CLK(clk),
    .D(_0961_),
    .RESET_B(net123),
    .Q(\mem[30][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9660_ (.CLK(clk),
    .D(_0962_),
    .RESET_B(net123),
    .Q(\mem[30][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9661_ (.CLK(clk),
    .D(_0963_),
    .RESET_B(net197),
    .Q(\mem[30][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9662_ (.CLK(clk),
    .D(_0964_),
    .RESET_B(net197),
    .Q(\mem[30][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9663_ (.CLK(clk),
    .D(_0965_),
    .RESET_B(net178),
    .Q(\mem[30][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9664_ (.CLK(clk),
    .D(_0966_),
    .RESET_B(net182),
    .Q(\mem[30][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9665_ (.CLK(clk),
    .D(_0967_),
    .RESET_B(net202),
    .Q(\mem[30][7] ));
 sky130_fd_sc_hd__dfrtp_1 _9666_ (.CLK(clk),
    .D(_0968_),
    .RESET_B(net201),
    .Q(\mem[30][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9667_ (.CLK(clk),
    .D(_0969_),
    .RESET_B(net203),
    .Q(\mem[30][9] ));
 sky130_fd_sc_hd__dfrtp_1 _9668_ (.CLK(clk),
    .D(_0970_),
    .RESET_B(net204),
    .Q(\mem[30][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9669_ (.CLK(clk),
    .D(_0971_),
    .RESET_B(net229),
    .Q(\mem[30][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9670_ (.CLK(clk),
    .D(_0972_),
    .RESET_B(net217),
    .Q(\mem[30][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9671_ (.CLK(clk),
    .D(_0973_),
    .RESET_B(net230),
    .Q(\mem[30][13] ));
 sky130_fd_sc_hd__dfrtp_1 _9672_ (.CLK(clk),
    .D(_0974_),
    .RESET_B(net232),
    .Q(\mem[30][14] ));
 sky130_fd_sc_hd__dfrtp_1 _9673_ (.CLK(clk),
    .D(_0975_),
    .RESET_B(net238),
    .Q(\mem[30][15] ));
 sky130_fd_sc_hd__dfrtp_1 _9674_ (.CLK(clk),
    .D(_0976_),
    .RESET_B(net232),
    .Q(\mem[30][16] ));
 sky130_fd_sc_hd__dfrtp_1 _9675_ (.CLK(clk),
    .D(_0977_),
    .RESET_B(net212),
    .Q(\mem[30][17] ));
 sky130_fd_sc_hd__dfrtp_1 _9676_ (.CLK(clk),
    .D(_0978_),
    .RESET_B(net162),
    .Q(\mem[30][18] ));
 sky130_fd_sc_hd__dfrtp_1 _9677_ (.CLK(clk),
    .D(_0979_),
    .RESET_B(net162),
    .Q(\mem[30][19] ));
 sky130_fd_sc_hd__dfrtp_1 _9678_ (.CLK(clk),
    .D(_0980_),
    .RESET_B(net165),
    .Q(\mem[30][20] ));
 sky130_fd_sc_hd__dfrtp_1 _9679_ (.CLK(clk),
    .D(_0981_),
    .RESET_B(net153),
    .Q(\mem[30][21] ));
 sky130_fd_sc_hd__dfrtp_1 _9680_ (.CLK(clk),
    .D(_0982_),
    .RESET_B(net146),
    .Q(\mem[30][22] ));
 sky130_fd_sc_hd__dfrtp_1 _9681_ (.CLK(clk),
    .D(_0983_),
    .RESET_B(net153),
    .Q(\mem[30][23] ));
 sky130_fd_sc_hd__dfrtp_1 _9682_ (.CLK(clk),
    .D(_0984_),
    .RESET_B(net153),
    .Q(\mem[30][24] ));
 sky130_fd_sc_hd__dfrtp_1 _9683_ (.CLK(clk),
    .D(_0985_),
    .RESET_B(net146),
    .Q(\mem[30][25] ));
 sky130_fd_sc_hd__dfrtp_1 _9684_ (.CLK(clk),
    .D(_0986_),
    .RESET_B(net144),
    .Q(\mem[30][26] ));
 sky130_fd_sc_hd__dfrtp_1 _9685_ (.CLK(clk),
    .D(_0987_),
    .RESET_B(net144),
    .Q(\mem[30][27] ));
 sky130_fd_sc_hd__dfrtp_1 _9686_ (.CLK(clk),
    .D(_0988_),
    .RESET_B(net119),
    .Q(\mem[30][28] ));
 sky130_fd_sc_hd__dfrtp_1 _9687_ (.CLK(clk),
    .D(_0989_),
    .RESET_B(net119),
    .Q(\mem[30][29] ));
 sky130_fd_sc_hd__dfrtp_1 _9688_ (.CLK(clk),
    .D(_0990_),
    .RESET_B(net116),
    .Q(\mem[30][30] ));
 sky130_fd_sc_hd__dfrtp_1 _9689_ (.CLK(clk),
    .D(_0991_),
    .RESET_B(net120),
    .Q(\mem[30][31] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14435 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(rd_addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(rd_addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(rd_addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_8 input4 (.A(rd_addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_8 input5 (.A(rd_addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(rd_addr1[0]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(rd_addr1[1]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(rd_addr1[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(rd_addr1[3]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(rd_addr1[4]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(we0),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(wr_addr0[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(wr_addr0[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(wr_addr0[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_6 input16 (.A(wr_addr0[3]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(wr_addr0[4]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(wr_din0[0]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(wr_din0[10]),
    .X(net19));
 sky130_fd_sc_hd__buf_8 input20 (.A(wr_din0[11]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_8 input21 (.A(wr_din0[12]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_16 input22 (.A(wr_din0[13]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(wr_din0[14]),
    .X(net23));
 sky130_fd_sc_hd__buf_6 input24 (.A(wr_din0[15]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(wr_din0[16]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(wr_din0[17]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(wr_din0[18]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_8 input28 (.A(wr_din0[19]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(wr_din0[1]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input30 (.A(wr_din0[20]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(wr_din0[21]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(wr_din0[22]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(wr_din0[23]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 input34 (.A(wr_din0[24]),
    .X(net34));
 sky130_fd_sc_hd__buf_8 input35 (.A(wr_din0[25]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(wr_din0[26]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(wr_din0[27]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(wr_din0[28]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(wr_din0[29]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input40 (.A(wr_din0[2]),
    .X(net40));
 sky130_fd_sc_hd__buf_4 input41 (.A(wr_din0[30]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(wr_din0[31]),
    .X(net42));
 sky130_fd_sc_hd__buf_6 input43 (.A(wr_din0[3]),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(wr_din0[4]),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(wr_din0[5]),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input46 (.A(wr_din0[6]),
    .X(net46));
 sky130_fd_sc_hd__buf_6 input47 (.A(wr_din0[7]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(wr_din0[8]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(wr_din0[9]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(rd_dout0[0]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(rd_dout0[10]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(rd_dout0[11]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(rd_dout0[12]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(rd_dout0[13]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(rd_dout0[14]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(rd_dout0[15]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(rd_dout0[16]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(rd_dout0[17]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(rd_dout0[18]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(rd_dout0[19]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(rd_dout0[1]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(rd_dout0[20]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(rd_dout0[21]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(rd_dout0[22]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(rd_dout0[23]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(rd_dout0[24]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(rd_dout0[25]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(rd_dout0[26]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(rd_dout0[27]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(rd_dout0[28]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(rd_dout0[29]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(rd_dout0[2]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(rd_dout0[30]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(rd_dout0[31]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(rd_dout0[3]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(rd_dout0[4]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(rd_dout0[5]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(rd_dout0[6]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(rd_dout0[7]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(rd_dout0[8]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(rd_dout0[9]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(rd_dout1[0]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(rd_dout1[10]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(rd_dout1[11]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(rd_dout1[12]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(rd_dout1[13]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(rd_dout1[14]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(rd_dout1[15]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(rd_dout1[16]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(rd_dout1[17]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(rd_dout1[18]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(rd_dout1[19]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(rd_dout1[1]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(rd_dout1[20]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(rd_dout1[21]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(rd_dout1[22]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(rd_dout1[23]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(rd_dout1[24]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(rd_dout1[25]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(rd_dout1[26]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(rd_dout1[27]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(rd_dout1[28]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(rd_dout1[29]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(rd_dout1[2]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(rd_dout1[30]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(rd_dout1[31]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(rd_dout1[3]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(rd_dout1[4]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(rd_dout1[5]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(rd_dout1[6]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(rd_dout1[7]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(rd_dout1[8]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(rd_dout1[9]));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(net121),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(net120),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(net120),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net120),
    .X(net118));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(net136),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net136),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net129),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net129),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net136),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net133),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net133),
    .X(net131));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net136),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net11),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 fanout139 (.A(net147),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net142),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 fanout142 (.A(net147),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net147),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 fanout144 (.A(net147),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(net147),
    .X(net145));
 sky130_fd_sc_hd__buf_2 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net173),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net151),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net173),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 fanout153 (.A(net173),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net156),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 fanout156 (.A(net173),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net164),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net164),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net164),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(net164),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net164),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net173),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net172),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 fanout168 (.A(net172),
    .X(net168));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(net172),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(net172),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net11),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net178),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_2 fanout178 (.A(net193),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 fanout181 (.A(net193),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net193),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 fanout183 (.A(net193),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(net192),
    .X(net184));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(net192),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net192),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net192),
    .X(net188));
 sky130_fd_sc_hd__buf_2 fanout189 (.A(net192),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net192),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net246),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net200),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net200),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net200),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net200),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_2 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net246),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net210),
    .X(net201));
 sky130_fd_sc_hd__buf_2 fanout202 (.A(net210),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net210),
    .X(net203));
 sky130_fd_sc_hd__buf_2 fanout204 (.A(net210),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net210),
    .X(net205));
 sky130_fd_sc_hd__buf_2 fanout206 (.A(net210),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net209),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(net246),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net213),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net218),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(net218),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net218),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout216 (.A(net218),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 fanout218 (.A(net228),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(net223),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net223),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(net228),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net228),
    .X(net224));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(net228),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_2 fanout228 (.A(net246),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net245),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(net245),
    .X(net231));
 sky130_fd_sc_hd__buf_2 fanout232 (.A(net245),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net237),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net237),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(net245),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net244),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_4 fanout240 (.A(net244),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net244),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 fanout242 (.A(net244),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_2 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net11),
    .X(net246));
endmodule
